*FIRST LINE IS A COMMENT

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.88 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u

.SUBCKT sram_rom_column_mux
+ bl bl_out sel gnd
* INOUT : bl 
* INOUT : bl_out 
* INOUT : sel 
* INOUT : gnd 
Xmux_tx1 bl sel bl_out gnd sky130_fd_pr__nfet_01v8 m=1 w=2.88 l=0.15 pd=6.06 ps=6.06 as=1.08u ad=1.08u
.ENDS sram_rom_column_mux

.SUBCKT sram_rom_column_mux_array
+ bl_0 bl_1 bl_2 bl_3 bl_4 bl_5 bl_6 bl_7 bl_8 bl_9 bl_10 bl_11 bl_12
+ bl_13 bl_14 bl_15 bl_16 bl_17 bl_18 bl_19 bl_20 bl_21 bl_22 bl_23
+ bl_24 bl_25 bl_26 bl_27 bl_28 bl_29 bl_30 bl_31 bl_32 bl_33 bl_34
+ bl_35 bl_36 bl_37 bl_38 bl_39 bl_40 bl_41 bl_42 bl_43 bl_44 bl_45
+ bl_46 bl_47 bl_48 bl_49 bl_50 bl_51 bl_52 bl_53 bl_54 bl_55 bl_56
+ bl_57 bl_58 bl_59 bl_60 bl_61 bl_62 bl_63 bl_64 bl_65 bl_66 bl_67
+ bl_68 bl_69 bl_70 bl_71 bl_72 bl_73 bl_74 bl_75 bl_76 bl_77 bl_78
+ bl_79 bl_80 bl_81 bl_82 bl_83 bl_84 bl_85 bl_86 bl_87 bl_88 bl_89
+ bl_90 bl_91 bl_92 bl_93 bl_94 bl_95 bl_96 bl_97 bl_98 bl_99 bl_100
+ bl_101 bl_102 bl_103 bl_104 bl_105 bl_106 bl_107 bl_108 bl_109 bl_110
+ bl_111 bl_112 bl_113 bl_114 bl_115 bl_116 bl_117 bl_118 bl_119 bl_120
+ bl_121 bl_122 bl_123 bl_124 bl_125 bl_126 bl_127 bl_128 bl_129 bl_130
+ bl_131 bl_132 bl_133 bl_134 bl_135 bl_136 bl_137 bl_138 bl_139 bl_140
+ bl_141 bl_142 bl_143 bl_144 bl_145 bl_146 bl_147 bl_148 bl_149 bl_150
+ bl_151 bl_152 bl_153 bl_154 bl_155 bl_156 bl_157 bl_158 bl_159 bl_160
+ bl_161 bl_162 bl_163 bl_164 bl_165 bl_166 bl_167 bl_168 bl_169 bl_170
+ bl_171 bl_172 bl_173 bl_174 bl_175 bl_176 bl_177 bl_178 bl_179 bl_180
+ bl_181 bl_182 bl_183 sel_0 sel_1 sel_2 sel_3 sel_4 sel_5 sel_6 sel_7
+ sel_8 sel_9 sel_10 sel_11 sel_12 sel_13 sel_14 sel_15 sel_16 sel_17
+ sel_18 sel_19 sel_20 sel_21 sel_22 bl_out_0 bl_out_1 bl_out_2 bl_out_3
+ bl_out_4 bl_out_5 bl_out_6 bl_out_7 gnd
* INOUT : bl_0 
* INOUT : bl_1 
* INOUT : bl_2 
* INOUT : bl_3 
* INOUT : bl_4 
* INOUT : bl_5 
* INOUT : bl_6 
* INOUT : bl_7 
* INOUT : bl_8 
* INOUT : bl_9 
* INOUT : bl_10 
* INOUT : bl_11 
* INOUT : bl_12 
* INOUT : bl_13 
* INOUT : bl_14 
* INOUT : bl_15 
* INOUT : bl_16 
* INOUT : bl_17 
* INOUT : bl_18 
* INOUT : bl_19 
* INOUT : bl_20 
* INOUT : bl_21 
* INOUT : bl_22 
* INOUT : bl_23 
* INOUT : bl_24 
* INOUT : bl_25 
* INOUT : bl_26 
* INOUT : bl_27 
* INOUT : bl_28 
* INOUT : bl_29 
* INOUT : bl_30 
* INOUT : bl_31 
* INOUT : bl_32 
* INOUT : bl_33 
* INOUT : bl_34 
* INOUT : bl_35 
* INOUT : bl_36 
* INOUT : bl_37 
* INOUT : bl_38 
* INOUT : bl_39 
* INOUT : bl_40 
* INOUT : bl_41 
* INOUT : bl_42 
* INOUT : bl_43 
* INOUT : bl_44 
* INOUT : bl_45 
* INOUT : bl_46 
* INOUT : bl_47 
* INOUT : bl_48 
* INOUT : bl_49 
* INOUT : bl_50 
* INOUT : bl_51 
* INOUT : bl_52 
* INOUT : bl_53 
* INOUT : bl_54 
* INOUT : bl_55 
* INOUT : bl_56 
* INOUT : bl_57 
* INOUT : bl_58 
* INOUT : bl_59 
* INOUT : bl_60 
* INOUT : bl_61 
* INOUT : bl_62 
* INOUT : bl_63 
* INOUT : bl_64 
* INOUT : bl_65 
* INOUT : bl_66 
* INOUT : bl_67 
* INOUT : bl_68 
* INOUT : bl_69 
* INOUT : bl_70 
* INOUT : bl_71 
* INOUT : bl_72 
* INOUT : bl_73 
* INOUT : bl_74 
* INOUT : bl_75 
* INOUT : bl_76 
* INOUT : bl_77 
* INOUT : bl_78 
* INOUT : bl_79 
* INOUT : bl_80 
* INOUT : bl_81 
* INOUT : bl_82 
* INOUT : bl_83 
* INOUT : bl_84 
* INOUT : bl_85 
* INOUT : bl_86 
* INOUT : bl_87 
* INOUT : bl_88 
* INOUT : bl_89 
* INOUT : bl_90 
* INOUT : bl_91 
* INOUT : bl_92 
* INOUT : bl_93 
* INOUT : bl_94 
* INOUT : bl_95 
* INOUT : bl_96 
* INOUT : bl_97 
* INOUT : bl_98 
* INOUT : bl_99 
* INOUT : bl_100 
* INOUT : bl_101 
* INOUT : bl_102 
* INOUT : bl_103 
* INOUT : bl_104 
* INOUT : bl_105 
* INOUT : bl_106 
* INOUT : bl_107 
* INOUT : bl_108 
* INOUT : bl_109 
* INOUT : bl_110 
* INOUT : bl_111 
* INOUT : bl_112 
* INOUT : bl_113 
* INOUT : bl_114 
* INOUT : bl_115 
* INOUT : bl_116 
* INOUT : bl_117 
* INOUT : bl_118 
* INOUT : bl_119 
* INOUT : bl_120 
* INOUT : bl_121 
* INOUT : bl_122 
* INOUT : bl_123 
* INOUT : bl_124 
* INOUT : bl_125 
* INOUT : bl_126 
* INOUT : bl_127 
* INOUT : bl_128 
* INOUT : bl_129 
* INOUT : bl_130 
* INOUT : bl_131 
* INOUT : bl_132 
* INOUT : bl_133 
* INOUT : bl_134 
* INOUT : bl_135 
* INOUT : bl_136 
* INOUT : bl_137 
* INOUT : bl_138 
* INOUT : bl_139 
* INOUT : bl_140 
* INOUT : bl_141 
* INOUT : bl_142 
* INOUT : bl_143 
* INOUT : bl_144 
* INOUT : bl_145 
* INOUT : bl_146 
* INOUT : bl_147 
* INOUT : bl_148 
* INOUT : bl_149 
* INOUT : bl_150 
* INOUT : bl_151 
* INOUT : bl_152 
* INOUT : bl_153 
* INOUT : bl_154 
* INOUT : bl_155 
* INOUT : bl_156 
* INOUT : bl_157 
* INOUT : bl_158 
* INOUT : bl_159 
* INOUT : bl_160 
* INOUT : bl_161 
* INOUT : bl_162 
* INOUT : bl_163 
* INOUT : bl_164 
* INOUT : bl_165 
* INOUT : bl_166 
* INOUT : bl_167 
* INOUT : bl_168 
* INOUT : bl_169 
* INOUT : bl_170 
* INOUT : bl_171 
* INOUT : bl_172 
* INOUT : bl_173 
* INOUT : bl_174 
* INOUT : bl_175 
* INOUT : bl_176 
* INOUT : bl_177 
* INOUT : bl_178 
* INOUT : bl_179 
* INOUT : bl_180 
* INOUT : bl_181 
* INOUT : bl_182 
* INOUT : bl_183 
* INOUT : sel_0 
* INOUT : sel_1 
* INOUT : sel_2 
* INOUT : sel_3 
* INOUT : sel_4 
* INOUT : sel_5 
* INOUT : sel_6 
* INOUT : sel_7 
* INOUT : sel_8 
* INOUT : sel_9 
* INOUT : sel_10 
* INOUT : sel_11 
* INOUT : sel_12 
* INOUT : sel_13 
* INOUT : sel_14 
* INOUT : sel_15 
* INOUT : sel_16 
* INOUT : sel_17 
* INOUT : sel_18 
* INOUT : sel_19 
* INOUT : sel_20 
* INOUT : sel_21 
* INOUT : sel_22 
* INOUT : bl_out_0 
* INOUT : bl_out_1 
* INOUT : bl_out_2 
* INOUT : bl_out_3 
* INOUT : bl_out_4 
* INOUT : bl_out_5 
* INOUT : bl_out_6 
* INOUT : bl_out_7 
* INOUT : gnd 
* cols: 184 word_size: 8 
XXMUX0
+ bl_0 bl_out_0 sel_0 gnd
+ sram_rom_column_mux
XXMUX1
+ bl_1 bl_out_0 sel_1 gnd
+ sram_rom_column_mux
XXMUX2
+ bl_2 bl_out_0 sel_2 gnd
+ sram_rom_column_mux
XXMUX3
+ bl_3 bl_out_0 sel_3 gnd
+ sram_rom_column_mux
XXMUX4
+ bl_4 bl_out_0 sel_4 gnd
+ sram_rom_column_mux
XXMUX5
+ bl_5 bl_out_0 sel_5 gnd
+ sram_rom_column_mux
XXMUX6
+ bl_6 bl_out_0 sel_6 gnd
+ sram_rom_column_mux
XXMUX7
+ bl_7 bl_out_0 sel_7 gnd
+ sram_rom_column_mux
XXMUX8
+ bl_8 bl_out_0 sel_8 gnd
+ sram_rom_column_mux
XXMUX9
+ bl_9 bl_out_0 sel_9 gnd
+ sram_rom_column_mux
XXMUX10
+ bl_10 bl_out_0 sel_10 gnd
+ sram_rom_column_mux
XXMUX11
+ bl_11 bl_out_0 sel_11 gnd
+ sram_rom_column_mux
XXMUX12
+ bl_12 bl_out_0 sel_12 gnd
+ sram_rom_column_mux
XXMUX13
+ bl_13 bl_out_0 sel_13 gnd
+ sram_rom_column_mux
XXMUX14
+ bl_14 bl_out_0 sel_14 gnd
+ sram_rom_column_mux
XXMUX15
+ bl_15 bl_out_0 sel_15 gnd
+ sram_rom_column_mux
XXMUX16
+ bl_16 bl_out_0 sel_16 gnd
+ sram_rom_column_mux
XXMUX17
+ bl_17 bl_out_0 sel_17 gnd
+ sram_rom_column_mux
XXMUX18
+ bl_18 bl_out_0 sel_18 gnd
+ sram_rom_column_mux
XXMUX19
+ bl_19 bl_out_0 sel_19 gnd
+ sram_rom_column_mux
XXMUX20
+ bl_20 bl_out_0 sel_20 gnd
+ sram_rom_column_mux
XXMUX21
+ bl_21 bl_out_0 sel_21 gnd
+ sram_rom_column_mux
XXMUX22
+ bl_22 bl_out_0 sel_22 gnd
+ sram_rom_column_mux
XXMUX23
+ bl_23 bl_out_1 sel_0 gnd
+ sram_rom_column_mux
XXMUX24
+ bl_24 bl_out_1 sel_1 gnd
+ sram_rom_column_mux
XXMUX25
+ bl_25 bl_out_1 sel_2 gnd
+ sram_rom_column_mux
XXMUX26
+ bl_26 bl_out_1 sel_3 gnd
+ sram_rom_column_mux
XXMUX27
+ bl_27 bl_out_1 sel_4 gnd
+ sram_rom_column_mux
XXMUX28
+ bl_28 bl_out_1 sel_5 gnd
+ sram_rom_column_mux
XXMUX29
+ bl_29 bl_out_1 sel_6 gnd
+ sram_rom_column_mux
XXMUX30
+ bl_30 bl_out_1 sel_7 gnd
+ sram_rom_column_mux
XXMUX31
+ bl_31 bl_out_1 sel_8 gnd
+ sram_rom_column_mux
XXMUX32
+ bl_32 bl_out_1 sel_9 gnd
+ sram_rom_column_mux
XXMUX33
+ bl_33 bl_out_1 sel_10 gnd
+ sram_rom_column_mux
XXMUX34
+ bl_34 bl_out_1 sel_11 gnd
+ sram_rom_column_mux
XXMUX35
+ bl_35 bl_out_1 sel_12 gnd
+ sram_rom_column_mux
XXMUX36
+ bl_36 bl_out_1 sel_13 gnd
+ sram_rom_column_mux
XXMUX37
+ bl_37 bl_out_1 sel_14 gnd
+ sram_rom_column_mux
XXMUX38
+ bl_38 bl_out_1 sel_15 gnd
+ sram_rom_column_mux
XXMUX39
+ bl_39 bl_out_1 sel_16 gnd
+ sram_rom_column_mux
XXMUX40
+ bl_40 bl_out_1 sel_17 gnd
+ sram_rom_column_mux
XXMUX41
+ bl_41 bl_out_1 sel_18 gnd
+ sram_rom_column_mux
XXMUX42
+ bl_42 bl_out_1 sel_19 gnd
+ sram_rom_column_mux
XXMUX43
+ bl_43 bl_out_1 sel_20 gnd
+ sram_rom_column_mux
XXMUX44
+ bl_44 bl_out_1 sel_21 gnd
+ sram_rom_column_mux
XXMUX45
+ bl_45 bl_out_1 sel_22 gnd
+ sram_rom_column_mux
XXMUX46
+ bl_46 bl_out_2 sel_0 gnd
+ sram_rom_column_mux
XXMUX47
+ bl_47 bl_out_2 sel_1 gnd
+ sram_rom_column_mux
XXMUX48
+ bl_48 bl_out_2 sel_2 gnd
+ sram_rom_column_mux
XXMUX49
+ bl_49 bl_out_2 sel_3 gnd
+ sram_rom_column_mux
XXMUX50
+ bl_50 bl_out_2 sel_4 gnd
+ sram_rom_column_mux
XXMUX51
+ bl_51 bl_out_2 sel_5 gnd
+ sram_rom_column_mux
XXMUX52
+ bl_52 bl_out_2 sel_6 gnd
+ sram_rom_column_mux
XXMUX53
+ bl_53 bl_out_2 sel_7 gnd
+ sram_rom_column_mux
XXMUX54
+ bl_54 bl_out_2 sel_8 gnd
+ sram_rom_column_mux
XXMUX55
+ bl_55 bl_out_2 sel_9 gnd
+ sram_rom_column_mux
XXMUX56
+ bl_56 bl_out_2 sel_10 gnd
+ sram_rom_column_mux
XXMUX57
+ bl_57 bl_out_2 sel_11 gnd
+ sram_rom_column_mux
XXMUX58
+ bl_58 bl_out_2 sel_12 gnd
+ sram_rom_column_mux
XXMUX59
+ bl_59 bl_out_2 sel_13 gnd
+ sram_rom_column_mux
XXMUX60
+ bl_60 bl_out_2 sel_14 gnd
+ sram_rom_column_mux
XXMUX61
+ bl_61 bl_out_2 sel_15 gnd
+ sram_rom_column_mux
XXMUX62
+ bl_62 bl_out_2 sel_16 gnd
+ sram_rom_column_mux
XXMUX63
+ bl_63 bl_out_2 sel_17 gnd
+ sram_rom_column_mux
XXMUX64
+ bl_64 bl_out_2 sel_18 gnd
+ sram_rom_column_mux
XXMUX65
+ bl_65 bl_out_2 sel_19 gnd
+ sram_rom_column_mux
XXMUX66
+ bl_66 bl_out_2 sel_20 gnd
+ sram_rom_column_mux
XXMUX67
+ bl_67 bl_out_2 sel_21 gnd
+ sram_rom_column_mux
XXMUX68
+ bl_68 bl_out_2 sel_22 gnd
+ sram_rom_column_mux
XXMUX69
+ bl_69 bl_out_3 sel_0 gnd
+ sram_rom_column_mux
XXMUX70
+ bl_70 bl_out_3 sel_1 gnd
+ sram_rom_column_mux
XXMUX71
+ bl_71 bl_out_3 sel_2 gnd
+ sram_rom_column_mux
XXMUX72
+ bl_72 bl_out_3 sel_3 gnd
+ sram_rom_column_mux
XXMUX73
+ bl_73 bl_out_3 sel_4 gnd
+ sram_rom_column_mux
XXMUX74
+ bl_74 bl_out_3 sel_5 gnd
+ sram_rom_column_mux
XXMUX75
+ bl_75 bl_out_3 sel_6 gnd
+ sram_rom_column_mux
XXMUX76
+ bl_76 bl_out_3 sel_7 gnd
+ sram_rom_column_mux
XXMUX77
+ bl_77 bl_out_3 sel_8 gnd
+ sram_rom_column_mux
XXMUX78
+ bl_78 bl_out_3 sel_9 gnd
+ sram_rom_column_mux
XXMUX79
+ bl_79 bl_out_3 sel_10 gnd
+ sram_rom_column_mux
XXMUX80
+ bl_80 bl_out_3 sel_11 gnd
+ sram_rom_column_mux
XXMUX81
+ bl_81 bl_out_3 sel_12 gnd
+ sram_rom_column_mux
XXMUX82
+ bl_82 bl_out_3 sel_13 gnd
+ sram_rom_column_mux
XXMUX83
+ bl_83 bl_out_3 sel_14 gnd
+ sram_rom_column_mux
XXMUX84
+ bl_84 bl_out_3 sel_15 gnd
+ sram_rom_column_mux
XXMUX85
+ bl_85 bl_out_3 sel_16 gnd
+ sram_rom_column_mux
XXMUX86
+ bl_86 bl_out_3 sel_17 gnd
+ sram_rom_column_mux
XXMUX87
+ bl_87 bl_out_3 sel_18 gnd
+ sram_rom_column_mux
XXMUX88
+ bl_88 bl_out_3 sel_19 gnd
+ sram_rom_column_mux
XXMUX89
+ bl_89 bl_out_3 sel_20 gnd
+ sram_rom_column_mux
XXMUX90
+ bl_90 bl_out_3 sel_21 gnd
+ sram_rom_column_mux
XXMUX91
+ bl_91 bl_out_3 sel_22 gnd
+ sram_rom_column_mux
XXMUX92
+ bl_92 bl_out_4 sel_0 gnd
+ sram_rom_column_mux
XXMUX93
+ bl_93 bl_out_4 sel_1 gnd
+ sram_rom_column_mux
XXMUX94
+ bl_94 bl_out_4 sel_2 gnd
+ sram_rom_column_mux
XXMUX95
+ bl_95 bl_out_4 sel_3 gnd
+ sram_rom_column_mux
XXMUX96
+ bl_96 bl_out_4 sel_4 gnd
+ sram_rom_column_mux
XXMUX97
+ bl_97 bl_out_4 sel_5 gnd
+ sram_rom_column_mux
XXMUX98
+ bl_98 bl_out_4 sel_6 gnd
+ sram_rom_column_mux
XXMUX99
+ bl_99 bl_out_4 sel_7 gnd
+ sram_rom_column_mux
XXMUX100
+ bl_100 bl_out_4 sel_8 gnd
+ sram_rom_column_mux
XXMUX101
+ bl_101 bl_out_4 sel_9 gnd
+ sram_rom_column_mux
XXMUX102
+ bl_102 bl_out_4 sel_10 gnd
+ sram_rom_column_mux
XXMUX103
+ bl_103 bl_out_4 sel_11 gnd
+ sram_rom_column_mux
XXMUX104
+ bl_104 bl_out_4 sel_12 gnd
+ sram_rom_column_mux
XXMUX105
+ bl_105 bl_out_4 sel_13 gnd
+ sram_rom_column_mux
XXMUX106
+ bl_106 bl_out_4 sel_14 gnd
+ sram_rom_column_mux
XXMUX107
+ bl_107 bl_out_4 sel_15 gnd
+ sram_rom_column_mux
XXMUX108
+ bl_108 bl_out_4 sel_16 gnd
+ sram_rom_column_mux
XXMUX109
+ bl_109 bl_out_4 sel_17 gnd
+ sram_rom_column_mux
XXMUX110
+ bl_110 bl_out_4 sel_18 gnd
+ sram_rom_column_mux
XXMUX111
+ bl_111 bl_out_4 sel_19 gnd
+ sram_rom_column_mux
XXMUX112
+ bl_112 bl_out_4 sel_20 gnd
+ sram_rom_column_mux
XXMUX113
+ bl_113 bl_out_4 sel_21 gnd
+ sram_rom_column_mux
XXMUX114
+ bl_114 bl_out_4 sel_22 gnd
+ sram_rom_column_mux
XXMUX115
+ bl_115 bl_out_5 sel_0 gnd
+ sram_rom_column_mux
XXMUX116
+ bl_116 bl_out_5 sel_1 gnd
+ sram_rom_column_mux
XXMUX117
+ bl_117 bl_out_5 sel_2 gnd
+ sram_rom_column_mux
XXMUX118
+ bl_118 bl_out_5 sel_3 gnd
+ sram_rom_column_mux
XXMUX119
+ bl_119 bl_out_5 sel_4 gnd
+ sram_rom_column_mux
XXMUX120
+ bl_120 bl_out_5 sel_5 gnd
+ sram_rom_column_mux
XXMUX121
+ bl_121 bl_out_5 sel_6 gnd
+ sram_rom_column_mux
XXMUX122
+ bl_122 bl_out_5 sel_7 gnd
+ sram_rom_column_mux
XXMUX123
+ bl_123 bl_out_5 sel_8 gnd
+ sram_rom_column_mux
XXMUX124
+ bl_124 bl_out_5 sel_9 gnd
+ sram_rom_column_mux
XXMUX125
+ bl_125 bl_out_5 sel_10 gnd
+ sram_rom_column_mux
XXMUX126
+ bl_126 bl_out_5 sel_11 gnd
+ sram_rom_column_mux
XXMUX127
+ bl_127 bl_out_5 sel_12 gnd
+ sram_rom_column_mux
XXMUX128
+ bl_128 bl_out_5 sel_13 gnd
+ sram_rom_column_mux
XXMUX129
+ bl_129 bl_out_5 sel_14 gnd
+ sram_rom_column_mux
XXMUX130
+ bl_130 bl_out_5 sel_15 gnd
+ sram_rom_column_mux
XXMUX131
+ bl_131 bl_out_5 sel_16 gnd
+ sram_rom_column_mux
XXMUX132
+ bl_132 bl_out_5 sel_17 gnd
+ sram_rom_column_mux
XXMUX133
+ bl_133 bl_out_5 sel_18 gnd
+ sram_rom_column_mux
XXMUX134
+ bl_134 bl_out_5 sel_19 gnd
+ sram_rom_column_mux
XXMUX135
+ bl_135 bl_out_5 sel_20 gnd
+ sram_rom_column_mux
XXMUX136
+ bl_136 bl_out_5 sel_21 gnd
+ sram_rom_column_mux
XXMUX137
+ bl_137 bl_out_5 sel_22 gnd
+ sram_rom_column_mux
XXMUX138
+ bl_138 bl_out_6 sel_0 gnd
+ sram_rom_column_mux
XXMUX139
+ bl_139 bl_out_6 sel_1 gnd
+ sram_rom_column_mux
XXMUX140
+ bl_140 bl_out_6 sel_2 gnd
+ sram_rom_column_mux
XXMUX141
+ bl_141 bl_out_6 sel_3 gnd
+ sram_rom_column_mux
XXMUX142
+ bl_142 bl_out_6 sel_4 gnd
+ sram_rom_column_mux
XXMUX143
+ bl_143 bl_out_6 sel_5 gnd
+ sram_rom_column_mux
XXMUX144
+ bl_144 bl_out_6 sel_6 gnd
+ sram_rom_column_mux
XXMUX145
+ bl_145 bl_out_6 sel_7 gnd
+ sram_rom_column_mux
XXMUX146
+ bl_146 bl_out_6 sel_8 gnd
+ sram_rom_column_mux
XXMUX147
+ bl_147 bl_out_6 sel_9 gnd
+ sram_rom_column_mux
XXMUX148
+ bl_148 bl_out_6 sel_10 gnd
+ sram_rom_column_mux
XXMUX149
+ bl_149 bl_out_6 sel_11 gnd
+ sram_rom_column_mux
XXMUX150
+ bl_150 bl_out_6 sel_12 gnd
+ sram_rom_column_mux
XXMUX151
+ bl_151 bl_out_6 sel_13 gnd
+ sram_rom_column_mux
XXMUX152
+ bl_152 bl_out_6 sel_14 gnd
+ sram_rom_column_mux
XXMUX153
+ bl_153 bl_out_6 sel_15 gnd
+ sram_rom_column_mux
XXMUX154
+ bl_154 bl_out_6 sel_16 gnd
+ sram_rom_column_mux
XXMUX155
+ bl_155 bl_out_6 sel_17 gnd
+ sram_rom_column_mux
XXMUX156
+ bl_156 bl_out_6 sel_18 gnd
+ sram_rom_column_mux
XXMUX157
+ bl_157 bl_out_6 sel_19 gnd
+ sram_rom_column_mux
XXMUX158
+ bl_158 bl_out_6 sel_20 gnd
+ sram_rom_column_mux
XXMUX159
+ bl_159 bl_out_6 sel_21 gnd
+ sram_rom_column_mux
XXMUX160
+ bl_160 bl_out_6 sel_22 gnd
+ sram_rom_column_mux
XXMUX161
+ bl_161 bl_out_7 sel_0 gnd
+ sram_rom_column_mux
XXMUX162
+ bl_162 bl_out_7 sel_1 gnd
+ sram_rom_column_mux
XXMUX163
+ bl_163 bl_out_7 sel_2 gnd
+ sram_rom_column_mux
XXMUX164
+ bl_164 bl_out_7 sel_3 gnd
+ sram_rom_column_mux
XXMUX165
+ bl_165 bl_out_7 sel_4 gnd
+ sram_rom_column_mux
XXMUX166
+ bl_166 bl_out_7 sel_5 gnd
+ sram_rom_column_mux
XXMUX167
+ bl_167 bl_out_7 sel_6 gnd
+ sram_rom_column_mux
XXMUX168
+ bl_168 bl_out_7 sel_7 gnd
+ sram_rom_column_mux
XXMUX169
+ bl_169 bl_out_7 sel_8 gnd
+ sram_rom_column_mux
XXMUX170
+ bl_170 bl_out_7 sel_9 gnd
+ sram_rom_column_mux
XXMUX171
+ bl_171 bl_out_7 sel_10 gnd
+ sram_rom_column_mux
XXMUX172
+ bl_172 bl_out_7 sel_11 gnd
+ sram_rom_column_mux
XXMUX173
+ bl_173 bl_out_7 sel_12 gnd
+ sram_rom_column_mux
XXMUX174
+ bl_174 bl_out_7 sel_13 gnd
+ sram_rom_column_mux
XXMUX175
+ bl_175 bl_out_7 sel_14 gnd
+ sram_rom_column_mux
XXMUX176
+ bl_176 bl_out_7 sel_15 gnd
+ sram_rom_column_mux
XXMUX177
+ bl_177 bl_out_7 sel_16 gnd
+ sram_rom_column_mux
XXMUX178
+ bl_178 bl_out_7 sel_17 gnd
+ sram_rom_column_mux
XXMUX179
+ bl_179 bl_out_7 sel_18 gnd
+ sram_rom_column_mux
XXMUX180
+ bl_180 bl_out_7 sel_19 gnd
+ sram_rom_column_mux
XXMUX181
+ bl_181 bl_out_7 sel_20 gnd
+ sram_rom_column_mux
XXMUX182
+ bl_182 bl_out_7 sel_21 gnd
+ sram_rom_column_mux
XXMUX183
+ bl_183 bl_out_7 sel_22 gnd
+ sram_rom_column_mux
.ENDS sram_rom_column_mux_array

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u

.SUBCKT sram_rom_base_one_cell
+ bl_h bl_l wl gnd
* INOUT : bl_h 
* INOUT : bl_l 
* INPUT : wl 
* GROUND: gnd 
Xsram_rom_base_one_cell_nmos bl_h wl bl_l gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS sram_rom_base_one_cell

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=0.42 l=0.15 pd=1.14 ps=1.14 as=0.16u ad=0.16u

.SUBCKT sram_precharge_cell
+ vdd gate bitline
* POWER : vdd 
* INPUT : gate 
* OUTPUT: bitline 
Xprecharge_pmos bitline gate vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=0.42 l=0.15 pd=1.14 ps=1.14 as=0.16u ad=0.16u
.ENDS sram_precharge_cell

.SUBCKT sram_rom_precharge_array_1
+ pre_bl0_out pre_bl1_out pre_bl2_out pre_bl3_out pre_bl4_out
+ pre_bl5_out pre_bl6_out pre_bl7_out pre_bl8_out pre_bl9_out
+ pre_bl10_out pre_bl11_out pre_bl12_out pre_bl13_out pre_bl14_out
+ pre_bl15_out pre_bl16_out pre_bl17_out pre_bl18_out pre_bl19_out
+ pre_bl20_out pre_bl21_out pre_bl22_out gate vdd
* OUTPUT: pre_bl0_out 
* OUTPUT: pre_bl1_out 
* OUTPUT: pre_bl2_out 
* OUTPUT: pre_bl3_out 
* OUTPUT: pre_bl4_out 
* OUTPUT: pre_bl5_out 
* OUTPUT: pre_bl6_out 
* OUTPUT: pre_bl7_out 
* OUTPUT: pre_bl8_out 
* OUTPUT: pre_bl9_out 
* OUTPUT: pre_bl10_out 
* OUTPUT: pre_bl11_out 
* OUTPUT: pre_bl12_out 
* OUTPUT: pre_bl13_out 
* OUTPUT: pre_bl14_out 
* OUTPUT: pre_bl15_out 
* OUTPUT: pre_bl16_out 
* OUTPUT: pre_bl17_out 
* OUTPUT: pre_bl18_out 
* OUTPUT: pre_bl19_out 
* OUTPUT: pre_bl20_out 
* OUTPUT: pre_bl21_out 
* OUTPUT: pre_bl22_out 
* INPUT : gate 
* POWER : vdd 
Xpmos_c0
+ vdd gate pre_bl0_out
+ sram_precharge_cell
Xpmos_c1
+ vdd gate pre_bl1_out
+ sram_precharge_cell
Xpmos_c2
+ vdd gate pre_bl2_out
+ sram_precharge_cell
Xpmos_c3
+ vdd gate pre_bl3_out
+ sram_precharge_cell
Xpmos_c4
+ vdd gate pre_bl4_out
+ sram_precharge_cell
Xpmos_c5
+ vdd gate pre_bl5_out
+ sram_precharge_cell
Xpmos_c6
+ vdd gate pre_bl6_out
+ sram_precharge_cell
Xpmos_c7
+ vdd gate pre_bl7_out
+ sram_precharge_cell
Xpmos_c8
+ vdd gate pre_bl8_out
+ sram_precharge_cell
Xpmos_c9
+ vdd gate pre_bl9_out
+ sram_precharge_cell
Xpmos_c10
+ vdd gate pre_bl10_out
+ sram_precharge_cell
Xpmos_c11
+ vdd gate pre_bl11_out
+ sram_precharge_cell
Xpmos_c12
+ vdd gate pre_bl12_out
+ sram_precharge_cell
Xpmos_c13
+ vdd gate pre_bl13_out
+ sram_precharge_cell
Xpmos_c14
+ vdd gate pre_bl14_out
+ sram_precharge_cell
Xpmos_c15
+ vdd gate pre_bl15_out
+ sram_precharge_cell
Xpmos_c16
+ vdd gate pre_bl16_out
+ sram_precharge_cell
Xpmos_c17
+ vdd gate pre_bl17_out
+ sram_precharge_cell
Xpmos_c18
+ vdd gate pre_bl18_out
+ sram_precharge_cell
Xpmos_c19
+ vdd gate pre_bl19_out
+ sram_precharge_cell
Xpmos_c20
+ vdd gate pre_bl20_out
+ sram_precharge_cell
Xpmos_c21
+ vdd gate pre_bl21_out
+ sram_precharge_cell
Xpmos_c22
+ vdd gate pre_bl22_out
+ sram_precharge_cell
.ENDS sram_rom_precharge_array_1

.SUBCKT sram_rom_base_zero_cell
+ bl wl gnd
* INOUT : bl 
* INPUT : wl 
* GROUND: gnd 
Xsram_rom_base_zero_cell_nmos bl wl bl gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS sram_rom_base_zero_cell

.SUBCKT sram_rom_column_decode_array
+ bl_0_0 bl_0_1 bl_0_2 bl_0_3 bl_0_4 bl_0_5 bl_0_6 bl_0_7 bl_0_8 bl_0_9
+ bl_0_10 bl_0_11 bl_0_12 bl_0_13 bl_0_14 bl_0_15 bl_0_16 bl_0_17
+ bl_0_18 bl_0_19 bl_0_20 bl_0_21 bl_0_22 wl_0_0 wl_0_1 wl_0_2 wl_0_3
+ wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 precharge vdd gnd
* OUTPUT: bl_0_0 
* OUTPUT: bl_0_1 
* OUTPUT: bl_0_2 
* OUTPUT: bl_0_3 
* OUTPUT: bl_0_4 
* OUTPUT: bl_0_5 
* OUTPUT: bl_0_6 
* OUTPUT: bl_0_7 
* OUTPUT: bl_0_8 
* OUTPUT: bl_0_9 
* OUTPUT: bl_0_10 
* OUTPUT: bl_0_11 
* OUTPUT: bl_0_12 
* OUTPUT: bl_0_13 
* OUTPUT: bl_0_14 
* OUTPUT: bl_0_15 
* OUTPUT: bl_0_16 
* OUTPUT: bl_0_17 
* OUTPUT: bl_0_18 
* OUTPUT: bl_0_19 
* OUTPUT: bl_0_20 
* OUTPUT: bl_0_21 
* OUTPUT: bl_0_22 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : precharge 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_int_0_0 bl_0_0 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c1
+ bl_int_0_1 bl_0_1 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c2
+ bl_int_0_2 bl_0_2 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c3
+ bl_int_0_3 bl_0_3 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c4
+ bl_int_0_4 bl_0_4 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c5
+ bl_int_0_5 bl_0_5 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c6
+ bl_int_0_6 bl_0_6 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c7
+ bl_int_0_7 bl_0_7 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c8
+ bl_int_0_8 bl_0_8 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c9
+ bl_int_0_9 bl_0_9 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c10
+ bl_int_0_10 bl_0_10 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c11
+ bl_int_0_11 bl_0_11 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c12
+ bl_int_0_12 bl_0_12 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c13
+ bl_int_0_13 bl_0_13 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c14
+ bl_int_0_14 bl_0_14 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c15
+ bl_int_0_15 bl_0_15 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c16
+ bl_0_16 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c17
+ bl_0_17 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c18
+ bl_0_18 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c19
+ bl_0_19 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c20
+ bl_0_20 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c21
+ bl_0_21 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c22
+ bl_0_22 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c0
+ bl_int_0_0 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c1
+ bl_int_0_1 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c2
+ bl_int_0_2 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c3
+ bl_int_0_3 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c4
+ bl_int_0_4 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c5
+ bl_int_0_5 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c6
+ bl_int_0_6 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c7
+ bl_int_0_7 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c8
+ bl_int_0_8 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c9
+ bl_int_0_9 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c10
+ bl_int_0_10 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c11
+ bl_int_0_11 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c12
+ bl_int_0_12 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c13
+ bl_int_0_13 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c14
+ bl_int_0_14 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c15
+ bl_int_0_15 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c16
+ bl_int_1_16 bl_0_16 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c17
+ bl_int_1_17 bl_0_17 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c18
+ bl_int_1_18 bl_0_18 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c19
+ bl_int_1_19 bl_0_19 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c20
+ bl_int_1_20 bl_0_20 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c21
+ bl_int_1_21 bl_0_21 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c22
+ bl_int_1_22 bl_0_22 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r2_c0
+ bl_int_2_0 bl_int_0_0 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c1
+ bl_int_2_1 bl_int_0_1 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c2
+ bl_int_2_2 bl_int_0_2 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c3
+ bl_int_2_3 bl_int_0_3 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c4
+ bl_int_2_4 bl_int_0_4 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c5
+ bl_int_2_5 bl_int_0_5 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c6
+ bl_int_2_6 bl_int_0_6 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c7
+ bl_int_2_7 bl_int_0_7 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c8
+ bl_int_0_8 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c9
+ bl_int_0_9 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c10
+ bl_int_0_10 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c11
+ bl_int_0_11 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c12
+ bl_int_0_12 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c13
+ bl_int_0_13 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c14
+ bl_int_0_14 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c15
+ bl_int_0_15 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c16
+ bl_int_2_16 bl_int_1_16 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c17
+ bl_int_2_17 bl_int_1_17 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c18
+ bl_int_2_18 bl_int_1_18 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c19
+ bl_int_2_19 bl_int_1_19 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c20
+ bl_int_2_20 bl_int_1_20 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c21
+ bl_int_2_21 bl_int_1_21 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c22
+ bl_int_2_22 bl_int_1_22 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r3_c0
+ bl_int_2_0 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c1
+ bl_int_2_1 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c2
+ bl_int_2_2 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c3
+ bl_int_2_3 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c4
+ bl_int_2_4 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c5
+ bl_int_2_5 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c6
+ bl_int_2_6 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c7
+ bl_int_2_7 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c8
+ bl_int_3_8 bl_int_0_8 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c9
+ bl_int_3_9 bl_int_0_9 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c10
+ bl_int_3_10 bl_int_0_10 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c11
+ bl_int_3_11 bl_int_0_11 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c12
+ bl_int_3_12 bl_int_0_12 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c13
+ bl_int_3_13 bl_int_0_13 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c14
+ bl_int_3_14 bl_int_0_14 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c15
+ bl_int_3_15 bl_int_0_15 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c16
+ bl_int_2_16 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c17
+ bl_int_2_17 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c18
+ bl_int_2_18 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c19
+ bl_int_2_19 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c20
+ bl_int_2_20 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c21
+ bl_int_2_21 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c22
+ bl_int_2_22 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c0
+ bl_int_4_0 bl_int_2_0 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c1
+ bl_int_4_1 bl_int_2_1 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c2
+ bl_int_4_2 bl_int_2_2 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c3
+ bl_int_4_3 bl_int_2_3 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c4
+ bl_int_2_4 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c5
+ bl_int_2_5 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c6
+ bl_int_2_6 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c7
+ bl_int_2_7 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c8
+ bl_int_4_8 bl_int_3_8 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c9
+ bl_int_4_9 bl_int_3_9 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c10
+ bl_int_4_10 bl_int_3_10 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c11
+ bl_int_4_11 bl_int_3_11 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c12
+ bl_int_3_12 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c13
+ bl_int_3_13 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c14
+ bl_int_3_14 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c15
+ bl_int_3_15 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c16
+ bl_int_4_16 bl_int_2_16 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c17
+ bl_int_4_17 bl_int_2_17 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c18
+ bl_int_4_18 bl_int_2_18 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c19
+ bl_int_4_19 bl_int_2_19 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c20
+ bl_int_2_20 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c21
+ bl_int_2_21 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c22
+ bl_int_2_22 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c0
+ bl_int_4_0 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c1
+ bl_int_4_1 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c2
+ bl_int_4_2 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c3
+ bl_int_4_3 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c4
+ bl_int_5_4 bl_int_2_4 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c5
+ bl_int_5_5 bl_int_2_5 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c6
+ bl_int_5_6 bl_int_2_6 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c7
+ bl_int_5_7 bl_int_2_7 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c8
+ bl_int_4_8 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c9
+ bl_int_4_9 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c10
+ bl_int_4_10 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c11
+ bl_int_4_11 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c12
+ bl_int_5_12 bl_int_3_12 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c13
+ bl_int_5_13 bl_int_3_13 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c14
+ bl_int_5_14 bl_int_3_14 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c15
+ bl_int_5_15 bl_int_3_15 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c16
+ bl_int_4_16 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c17
+ bl_int_4_17 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c18
+ bl_int_4_18 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c19
+ bl_int_4_19 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c20
+ bl_int_5_20 bl_int_2_20 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c21
+ bl_int_5_21 bl_int_2_21 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c22
+ bl_int_5_22 bl_int_2_22 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r6_c0
+ bl_int_6_0 bl_int_4_0 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c1
+ bl_int_6_1 bl_int_4_1 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c2
+ bl_int_4_2 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c3
+ bl_int_4_3 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c4
+ bl_int_6_4 bl_int_5_4 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c5
+ bl_int_6_5 bl_int_5_5 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c6
+ bl_int_5_6 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c7
+ bl_int_5_7 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c8
+ bl_int_6_8 bl_int_4_8 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c9
+ bl_int_6_9 bl_int_4_9 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c10
+ bl_int_4_10 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c11
+ bl_int_4_11 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c12
+ bl_int_6_12 bl_int_5_12 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c13
+ bl_int_6_13 bl_int_5_13 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c14
+ bl_int_5_14 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c15
+ bl_int_5_15 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c16
+ bl_int_6_16 bl_int_4_16 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c17
+ bl_int_6_17 bl_int_4_17 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c18
+ bl_int_4_18 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c19
+ bl_int_4_19 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c20
+ bl_int_6_20 bl_int_5_20 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c21
+ bl_int_6_21 bl_int_5_21 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c22
+ bl_int_5_22 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c0
+ bl_int_6_0 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c1
+ bl_int_6_1 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c2
+ bl_int_7_2 bl_int_4_2 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c3
+ bl_int_7_3 bl_int_4_3 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c4
+ bl_int_6_4 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c5
+ bl_int_6_5 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c6
+ bl_int_7_6 bl_int_5_6 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c7
+ bl_int_7_7 bl_int_5_7 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c8
+ bl_int_6_8 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c9
+ bl_int_6_9 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c10
+ bl_int_7_10 bl_int_4_10 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c11
+ bl_int_7_11 bl_int_4_11 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c12
+ bl_int_6_12 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c13
+ bl_int_6_13 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c14
+ bl_int_7_14 bl_int_5_14 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c15
+ bl_int_7_15 bl_int_5_15 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c16
+ bl_int_6_16 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c17
+ bl_int_6_17 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c18
+ bl_int_7_18 bl_int_4_18 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c19
+ bl_int_7_19 bl_int_4_19 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c20
+ bl_int_6_20 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c21
+ bl_int_6_21 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c22
+ bl_int_7_22 bl_int_5_22 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r8_c0
+ bl_int_8_0 bl_int_6_0 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c1
+ bl_int_6_1 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c2
+ bl_int_8_2 bl_int_7_2 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c3
+ bl_int_7_3 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c4
+ bl_int_8_4 bl_int_6_4 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c5
+ bl_int_6_5 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c6
+ bl_int_8_6 bl_int_7_6 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c7
+ bl_int_7_7 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c8
+ bl_int_8_8 bl_int_6_8 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c9
+ bl_int_6_9 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c10
+ bl_int_8_10 bl_int_7_10 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c11
+ bl_int_7_11 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c12
+ bl_int_8_12 bl_int_6_12 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c13
+ bl_int_6_13 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c14
+ bl_int_8_14 bl_int_7_14 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c15
+ bl_int_7_15 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c16
+ bl_int_8_16 bl_int_6_16 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c17
+ bl_int_6_17 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c18
+ bl_int_8_18 bl_int_7_18 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c19
+ bl_int_7_19 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c20
+ bl_int_8_20 bl_int_6_20 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c21
+ bl_int_6_21 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c22
+ bl_int_8_22 bl_int_7_22 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r9_c0
+ bl_int_8_0 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c1
+ bl_int_9_1 bl_int_6_1 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c2
+ bl_int_8_2 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c3
+ bl_int_9_3 bl_int_7_3 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c4
+ bl_int_8_4 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c5
+ bl_int_9_5 bl_int_6_5 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c6
+ bl_int_8_6 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c7
+ bl_int_9_7 bl_int_7_7 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c8
+ bl_int_8_8 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c9
+ bl_int_9_9 bl_int_6_9 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c10
+ bl_int_8_10 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c11
+ bl_int_9_11 bl_int_7_11 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c12
+ bl_int_8_12 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c13
+ bl_int_9_13 bl_int_6_13 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c14
+ bl_int_8_14 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c15
+ bl_int_9_15 bl_int_7_15 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c16
+ bl_int_8_16 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c17
+ bl_int_9_17 bl_int_6_17 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c18
+ bl_int_8_18 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c19
+ bl_int_9_19 bl_int_7_19 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c20
+ bl_int_8_20 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c21
+ bl_int_9_21 bl_int_6_21 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c22
+ bl_int_8_22 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c0
+ gnd bl_int_8_0 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c1
+ gnd bl_int_9_1 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c2
+ gnd bl_int_8_2 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c3
+ gnd bl_int_9_3 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c4
+ gnd bl_int_8_4 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c5
+ gnd bl_int_9_5 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c6
+ gnd bl_int_8_6 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c7
+ gnd bl_int_9_7 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c8
+ gnd bl_int_8_8 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c9
+ gnd bl_int_9_9 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c10
+ gnd bl_int_8_10 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c11
+ gnd bl_int_9_11 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c12
+ gnd bl_int_8_12 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c13
+ gnd bl_int_9_13 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c14
+ gnd bl_int_8_14 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c15
+ gnd bl_int_9_15 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c16
+ gnd bl_int_8_16 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c17
+ gnd bl_int_9_17 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c18
+ gnd bl_int_8_18 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c19
+ gnd bl_int_9_19 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c20
+ gnd bl_int_8_20 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c21
+ gnd bl_int_9_21 precharge gnd
+ sram_rom_base_one_cell
Xbit_r10_c22
+ gnd bl_int_8_22 precharge gnd
+ sram_rom_base_one_cell
Xbitcell_array_precharge
+ bl_0_0 bl_0_1 bl_0_2 bl_0_3 bl_0_4 bl_0_5 bl_0_6 bl_0_7 bl_0_8 bl_0_9
+ bl_0_10 bl_0_11 bl_0_12 bl_0_13 bl_0_14 bl_0_15 bl_0_16 bl_0_17
+ bl_0_18 bl_0_19 bl_0_20 bl_0_21 bl_0_22 precharge vdd
+ sram_rom_precharge_array_1
.ENDS sram_rom_column_decode_array
* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

* NGSPICE file created from sky130_fd_bd_sram__openram_sp_nand2_dec.ext - technology: EFS8A


* Top level circuit sky130_fd_bd_sram__openram_sp_nand2_dec
.subckt sky130_fd_bd_sram__openram_sp_nand2_dec A B Z VDD GND

X1001 Z B VDD VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1002 VDD A Z VDD sky130_fd_pr__pfet_01v8 W=1.12 L=0.15
X1000 Z A a_n722_276# GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
X1003 a_n722_276# B GND GND sky130_fd_pr__nfet_01v8 W=0.74 L=0.15
.ends


* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

.SUBCKT sram_inv_array_mod
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u
.ENDS sram_inv_array_mod

.SUBCKT sram_rom_address_control_buf
+ A_in A_out Abar_out clk vdd gnd
* INPUT : A_in 
* INOUT : A_out 
* OUTPUT: Abar_out 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
XXinvAbar
+ A_in Abar_internal vdd gnd
+ sram_inv_array_mod
XXnand_addr
+ clk Abar_internal A_out vdd gnd
+ sky130_fd_bd_sram__openram_sp_nand2_dec
XXnand_addr_bar
+ clk A_out Abar_out vdd gnd
+ sky130_fd_bd_sram__openram_sp_nand2_dec
.ENDS sram_rom_address_control_buf

.SUBCKT sram_rom_address_control_array_0
+ A0_in A1_in A2_in A3_in A4_in A0_out A1_out A2_out A3_out A4_out
+ Abar0_out Abar1_out Abar2_out Abar3_out Abar4_out clk vdd gnd
* INPUT : A0_in 
* INPUT : A1_in 
* INPUT : A2_in 
* INPUT : A3_in 
* INPUT : A4_in 
* OUTPUT: A0_out 
* OUTPUT: A1_out 
* OUTPUT: A2_out 
* OUTPUT: A3_out 
* OUTPUT: A4_out 
* OUTPUT: Abar0_out 
* OUTPUT: Abar1_out 
* OUTPUT: Abar2_out 
* OUTPUT: Abar3_out 
* OUTPUT: Abar4_out 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
XXaddr_buf_0
+ A0_in A0_out Abar0_out clk vdd gnd
+ sram_rom_address_control_buf
XXaddr_buf_1
+ A1_in A1_out Abar1_out clk vdd gnd
+ sram_rom_address_control_buf
XXaddr_buf_2
+ A2_in A2_out Abar2_out clk vdd gnd
+ sram_rom_address_control_buf
XXaddr_buf_3
+ A3_in A3_out Abar3_out clk vdd gnd
+ sram_rom_address_control_buf
XXaddr_buf_4
+ A4_in A4_out Abar4_out clk vdd gnd
+ sram_rom_address_control_buf
.ENDS sram_rom_address_control_array_0

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u

.SUBCKT sram_pinv_dec_2
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS sram_pinv_dec_2

.SUBCKT sram_rom_column_decode_wordline_buffer
+ in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12
+ in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 out_0
+ out_1 out_2 out_3 out_4 out_5 out_6 out_7 out_8 out_9 out_10 out_11
+ out_12 out_13 out_14 out_15 out_16 out_17 out_18 out_19 out_20 out_21
+ out_22 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* OUTPUT: out_8 
* OUTPUT: out_9 
* OUTPUT: out_10 
* OUTPUT: out_11 
* OUTPUT: out_12 
* OUTPUT: out_13 
* OUTPUT: out_14 
* OUTPUT: out_15 
* OUTPUT: out_16 
* OUTPUT: out_17 
* OUTPUT: out_18 
* OUTPUT: out_19 
* OUTPUT: out_20 
* OUTPUT: out_21 
* OUTPUT: out_22 
* POWER : vdd 
* GROUND: gnd 
* rows: 23 Buffer size of: 2
Xwld0
+ in_0 out_0 vdd gnd
+ sram_pinv_dec_2
Xwld1
+ in_1 out_1 vdd gnd
+ sram_pinv_dec_2
Xwld2
+ in_2 out_2 vdd gnd
+ sram_pinv_dec_2
Xwld3
+ in_3 out_3 vdd gnd
+ sram_pinv_dec_2
Xwld4
+ in_4 out_4 vdd gnd
+ sram_pinv_dec_2
Xwld5
+ in_5 out_5 vdd gnd
+ sram_pinv_dec_2
Xwld6
+ in_6 out_6 vdd gnd
+ sram_pinv_dec_2
Xwld7
+ in_7 out_7 vdd gnd
+ sram_pinv_dec_2
Xwld8
+ in_8 out_8 vdd gnd
+ sram_pinv_dec_2
Xwld9
+ in_9 out_9 vdd gnd
+ sram_pinv_dec_2
Xwld10
+ in_10 out_10 vdd gnd
+ sram_pinv_dec_2
Xwld11
+ in_11 out_11 vdd gnd
+ sram_pinv_dec_2
Xwld12
+ in_12 out_12 vdd gnd
+ sram_pinv_dec_2
Xwld13
+ in_13 out_13 vdd gnd
+ sram_pinv_dec_2
Xwld14
+ in_14 out_14 vdd gnd
+ sram_pinv_dec_2
Xwld15
+ in_15 out_15 vdd gnd
+ sram_pinv_dec_2
Xwld16
+ in_16 out_16 vdd gnd
+ sram_pinv_dec_2
Xwld17
+ in_17 out_17 vdd gnd
+ sram_pinv_dec_2
Xwld18
+ in_18 out_18 vdd gnd
+ sram_pinv_dec_2
Xwld19
+ in_19 out_19 vdd gnd
+ sram_pinv_dec_2
Xwld20
+ in_20 out_20 vdd gnd
+ sram_pinv_dec_2
Xwld21
+ in_21 out_21 vdd gnd
+ sram_pinv_dec_2
Xwld22
+ in_22 out_22 vdd gnd
+ sram_pinv_dec_2
.ENDS sram_rom_column_decode_wordline_buffer

.SUBCKT sram_rom_column_decode
+ A0 A1 A2 A3 A4 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10
+ wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21
+ wl_22 precharge clk vdd gnd
* INPUT : A0 
* INPUT : A1 
* INPUT : A2 
* INPUT : A3 
* INPUT : A4 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* INPUT : precharge 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
Xdecode_array_inst
+ wl_int0 wl_int1 wl_int2 wl_int3 wl_int4 wl_int5 wl_int6 wl_int7
+ wl_int8 wl_int9 wl_int10 wl_int11 wl_int12 wl_int13 wl_int14 wl_int15
+ wl_int16 wl_int17 wl_int18 wl_int19 wl_int20 wl_int21 wl_int22
+ Ab_int_4 A_int_4 Ab_int_3 A_int_3 Ab_int_2 A_int_2 Ab_int_1 A_int_1
+ Ab_int_0 A_int_0 precharge vdd gnd
+ sram_rom_column_decode_array
Xpre_control_array
+ A0 A1 A2 A3 A4 A_int_0 A_int_1 A_int_2 A_int_3 A_int_4 Ab_int_0
+ Ab_int_1 Ab_int_2 Ab_int_3 Ab_int_4 clk vdd gnd
+ sram_rom_address_control_array_0
Xrom_wordline_driver
+ wl_int0 wl_int1 wl_int2 wl_int3 wl_int4 wl_int5 wl_int6 wl_int7
+ wl_int8 wl_int9 wl_int10 wl_int11 wl_int12 wl_int13 wl_int14 wl_int15
+ wl_int16 wl_int17 wl_int18 wl_int19 wl_int20 wl_int21 wl_int22 wl_0
+ wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13
+ wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 vdd gnd
+ sram_rom_column_decode_wordline_buffer
.ENDS sram_rom_column_decode

.SUBCKT sram_pinv_dec_3
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u
.ENDS sram_pinv_dec_3

.SUBCKT sram_rom_bitline_inverter
+ in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12
+ in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 in_23
+ in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34
+ in_35 in_36 in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45
+ in_46 in_47 in_48 in_49 in_50 in_51 in_52 in_53 in_54 in_55 in_56
+ in_57 in_58 in_59 in_60 in_61 in_62 in_63 in_64 in_65 in_66 in_67
+ in_68 in_69 in_70 in_71 in_72 in_73 in_74 in_75 in_76 in_77 in_78
+ in_79 in_80 in_81 in_82 in_83 in_84 in_85 in_86 in_87 in_88 in_89
+ in_90 in_91 in_92 in_93 in_94 in_95 in_96 in_97 in_98 in_99 in_100
+ in_101 in_102 in_103 in_104 in_105 in_106 in_107 in_108 in_109 in_110
+ in_111 in_112 in_113 in_114 in_115 in_116 in_117 in_118 in_119 in_120
+ in_121 in_122 in_123 in_124 in_125 in_126 in_127 in_128 in_129 in_130
+ in_131 in_132 in_133 in_134 in_135 in_136 in_137 in_138 in_139 in_140
+ in_141 in_142 in_143 in_144 in_145 in_146 in_147 in_148 in_149 in_150
+ in_151 in_152 in_153 in_154 in_155 in_156 in_157 in_158 in_159 in_160
+ in_161 in_162 in_163 in_164 in_165 in_166 in_167 in_168 in_169 in_170
+ in_171 in_172 in_173 in_174 in_175 in_176 in_177 in_178 in_179 in_180
+ in_181 in_182 in_183 out_0 out_1 out_2 out_3 out_4 out_5 out_6 out_7
+ out_8 out_9 out_10 out_11 out_12 out_13 out_14 out_15 out_16 out_17
+ out_18 out_19 out_20 out_21 out_22 out_23 out_24 out_25 out_26 out_27
+ out_28 out_29 out_30 out_31 out_32 out_33 out_34 out_35 out_36 out_37
+ out_38 out_39 out_40 out_41 out_42 out_43 out_44 out_45 out_46 out_47
+ out_48 out_49 out_50 out_51 out_52 out_53 out_54 out_55 out_56 out_57
+ out_58 out_59 out_60 out_61 out_62 out_63 out_64 out_65 out_66 out_67
+ out_68 out_69 out_70 out_71 out_72 out_73 out_74 out_75 out_76 out_77
+ out_78 out_79 out_80 out_81 out_82 out_83 out_84 out_85 out_86 out_87
+ out_88 out_89 out_90 out_91 out_92 out_93 out_94 out_95 out_96 out_97
+ out_98 out_99 out_100 out_101 out_102 out_103 out_104 out_105 out_106
+ out_107 out_108 out_109 out_110 out_111 out_112 out_113 out_114
+ out_115 out_116 out_117 out_118 out_119 out_120 out_121 out_122
+ out_123 out_124 out_125 out_126 out_127 out_128 out_129 out_130
+ out_131 out_132 out_133 out_134 out_135 out_136 out_137 out_138
+ out_139 out_140 out_141 out_142 out_143 out_144 out_145 out_146
+ out_147 out_148 out_149 out_150 out_151 out_152 out_153 out_154
+ out_155 out_156 out_157 out_158 out_159 out_160 out_161 out_162
+ out_163 out_164 out_165 out_166 out_167 out_168 out_169 out_170
+ out_171 out_172 out_173 out_174 out_175 out_176 out_177 out_178
+ out_179 out_180 out_181 out_182 out_183 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* INPUT : in_23 
* INPUT : in_24 
* INPUT : in_25 
* INPUT : in_26 
* INPUT : in_27 
* INPUT : in_28 
* INPUT : in_29 
* INPUT : in_30 
* INPUT : in_31 
* INPUT : in_32 
* INPUT : in_33 
* INPUT : in_34 
* INPUT : in_35 
* INPUT : in_36 
* INPUT : in_37 
* INPUT : in_38 
* INPUT : in_39 
* INPUT : in_40 
* INPUT : in_41 
* INPUT : in_42 
* INPUT : in_43 
* INPUT : in_44 
* INPUT : in_45 
* INPUT : in_46 
* INPUT : in_47 
* INPUT : in_48 
* INPUT : in_49 
* INPUT : in_50 
* INPUT : in_51 
* INPUT : in_52 
* INPUT : in_53 
* INPUT : in_54 
* INPUT : in_55 
* INPUT : in_56 
* INPUT : in_57 
* INPUT : in_58 
* INPUT : in_59 
* INPUT : in_60 
* INPUT : in_61 
* INPUT : in_62 
* INPUT : in_63 
* INPUT : in_64 
* INPUT : in_65 
* INPUT : in_66 
* INPUT : in_67 
* INPUT : in_68 
* INPUT : in_69 
* INPUT : in_70 
* INPUT : in_71 
* INPUT : in_72 
* INPUT : in_73 
* INPUT : in_74 
* INPUT : in_75 
* INPUT : in_76 
* INPUT : in_77 
* INPUT : in_78 
* INPUT : in_79 
* INPUT : in_80 
* INPUT : in_81 
* INPUT : in_82 
* INPUT : in_83 
* INPUT : in_84 
* INPUT : in_85 
* INPUT : in_86 
* INPUT : in_87 
* INPUT : in_88 
* INPUT : in_89 
* INPUT : in_90 
* INPUT : in_91 
* INPUT : in_92 
* INPUT : in_93 
* INPUT : in_94 
* INPUT : in_95 
* INPUT : in_96 
* INPUT : in_97 
* INPUT : in_98 
* INPUT : in_99 
* INPUT : in_100 
* INPUT : in_101 
* INPUT : in_102 
* INPUT : in_103 
* INPUT : in_104 
* INPUT : in_105 
* INPUT : in_106 
* INPUT : in_107 
* INPUT : in_108 
* INPUT : in_109 
* INPUT : in_110 
* INPUT : in_111 
* INPUT : in_112 
* INPUT : in_113 
* INPUT : in_114 
* INPUT : in_115 
* INPUT : in_116 
* INPUT : in_117 
* INPUT : in_118 
* INPUT : in_119 
* INPUT : in_120 
* INPUT : in_121 
* INPUT : in_122 
* INPUT : in_123 
* INPUT : in_124 
* INPUT : in_125 
* INPUT : in_126 
* INPUT : in_127 
* INPUT : in_128 
* INPUT : in_129 
* INPUT : in_130 
* INPUT : in_131 
* INPUT : in_132 
* INPUT : in_133 
* INPUT : in_134 
* INPUT : in_135 
* INPUT : in_136 
* INPUT : in_137 
* INPUT : in_138 
* INPUT : in_139 
* INPUT : in_140 
* INPUT : in_141 
* INPUT : in_142 
* INPUT : in_143 
* INPUT : in_144 
* INPUT : in_145 
* INPUT : in_146 
* INPUT : in_147 
* INPUT : in_148 
* INPUT : in_149 
* INPUT : in_150 
* INPUT : in_151 
* INPUT : in_152 
* INPUT : in_153 
* INPUT : in_154 
* INPUT : in_155 
* INPUT : in_156 
* INPUT : in_157 
* INPUT : in_158 
* INPUT : in_159 
* INPUT : in_160 
* INPUT : in_161 
* INPUT : in_162 
* INPUT : in_163 
* INPUT : in_164 
* INPUT : in_165 
* INPUT : in_166 
* INPUT : in_167 
* INPUT : in_168 
* INPUT : in_169 
* INPUT : in_170 
* INPUT : in_171 
* INPUT : in_172 
* INPUT : in_173 
* INPUT : in_174 
* INPUT : in_175 
* INPUT : in_176 
* INPUT : in_177 
* INPUT : in_178 
* INPUT : in_179 
* INPUT : in_180 
* INPUT : in_181 
* INPUT : in_182 
* INPUT : in_183 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* OUTPUT: out_8 
* OUTPUT: out_9 
* OUTPUT: out_10 
* OUTPUT: out_11 
* OUTPUT: out_12 
* OUTPUT: out_13 
* OUTPUT: out_14 
* OUTPUT: out_15 
* OUTPUT: out_16 
* OUTPUT: out_17 
* OUTPUT: out_18 
* OUTPUT: out_19 
* OUTPUT: out_20 
* OUTPUT: out_21 
* OUTPUT: out_22 
* OUTPUT: out_23 
* OUTPUT: out_24 
* OUTPUT: out_25 
* OUTPUT: out_26 
* OUTPUT: out_27 
* OUTPUT: out_28 
* OUTPUT: out_29 
* OUTPUT: out_30 
* OUTPUT: out_31 
* OUTPUT: out_32 
* OUTPUT: out_33 
* OUTPUT: out_34 
* OUTPUT: out_35 
* OUTPUT: out_36 
* OUTPUT: out_37 
* OUTPUT: out_38 
* OUTPUT: out_39 
* OUTPUT: out_40 
* OUTPUT: out_41 
* OUTPUT: out_42 
* OUTPUT: out_43 
* OUTPUT: out_44 
* OUTPUT: out_45 
* OUTPUT: out_46 
* OUTPUT: out_47 
* OUTPUT: out_48 
* OUTPUT: out_49 
* OUTPUT: out_50 
* OUTPUT: out_51 
* OUTPUT: out_52 
* OUTPUT: out_53 
* OUTPUT: out_54 
* OUTPUT: out_55 
* OUTPUT: out_56 
* OUTPUT: out_57 
* OUTPUT: out_58 
* OUTPUT: out_59 
* OUTPUT: out_60 
* OUTPUT: out_61 
* OUTPUT: out_62 
* OUTPUT: out_63 
* OUTPUT: out_64 
* OUTPUT: out_65 
* OUTPUT: out_66 
* OUTPUT: out_67 
* OUTPUT: out_68 
* OUTPUT: out_69 
* OUTPUT: out_70 
* OUTPUT: out_71 
* OUTPUT: out_72 
* OUTPUT: out_73 
* OUTPUT: out_74 
* OUTPUT: out_75 
* OUTPUT: out_76 
* OUTPUT: out_77 
* OUTPUT: out_78 
* OUTPUT: out_79 
* OUTPUT: out_80 
* OUTPUT: out_81 
* OUTPUT: out_82 
* OUTPUT: out_83 
* OUTPUT: out_84 
* OUTPUT: out_85 
* OUTPUT: out_86 
* OUTPUT: out_87 
* OUTPUT: out_88 
* OUTPUT: out_89 
* OUTPUT: out_90 
* OUTPUT: out_91 
* OUTPUT: out_92 
* OUTPUT: out_93 
* OUTPUT: out_94 
* OUTPUT: out_95 
* OUTPUT: out_96 
* OUTPUT: out_97 
* OUTPUT: out_98 
* OUTPUT: out_99 
* OUTPUT: out_100 
* OUTPUT: out_101 
* OUTPUT: out_102 
* OUTPUT: out_103 
* OUTPUT: out_104 
* OUTPUT: out_105 
* OUTPUT: out_106 
* OUTPUT: out_107 
* OUTPUT: out_108 
* OUTPUT: out_109 
* OUTPUT: out_110 
* OUTPUT: out_111 
* OUTPUT: out_112 
* OUTPUT: out_113 
* OUTPUT: out_114 
* OUTPUT: out_115 
* OUTPUT: out_116 
* OUTPUT: out_117 
* OUTPUT: out_118 
* OUTPUT: out_119 
* OUTPUT: out_120 
* OUTPUT: out_121 
* OUTPUT: out_122 
* OUTPUT: out_123 
* OUTPUT: out_124 
* OUTPUT: out_125 
* OUTPUT: out_126 
* OUTPUT: out_127 
* OUTPUT: out_128 
* OUTPUT: out_129 
* OUTPUT: out_130 
* OUTPUT: out_131 
* OUTPUT: out_132 
* OUTPUT: out_133 
* OUTPUT: out_134 
* OUTPUT: out_135 
* OUTPUT: out_136 
* OUTPUT: out_137 
* OUTPUT: out_138 
* OUTPUT: out_139 
* OUTPUT: out_140 
* OUTPUT: out_141 
* OUTPUT: out_142 
* OUTPUT: out_143 
* OUTPUT: out_144 
* OUTPUT: out_145 
* OUTPUT: out_146 
* OUTPUT: out_147 
* OUTPUT: out_148 
* OUTPUT: out_149 
* OUTPUT: out_150 
* OUTPUT: out_151 
* OUTPUT: out_152 
* OUTPUT: out_153 
* OUTPUT: out_154 
* OUTPUT: out_155 
* OUTPUT: out_156 
* OUTPUT: out_157 
* OUTPUT: out_158 
* OUTPUT: out_159 
* OUTPUT: out_160 
* OUTPUT: out_161 
* OUTPUT: out_162 
* OUTPUT: out_163 
* OUTPUT: out_164 
* OUTPUT: out_165 
* OUTPUT: out_166 
* OUTPUT: out_167 
* OUTPUT: out_168 
* OUTPUT: out_169 
* OUTPUT: out_170 
* OUTPUT: out_171 
* OUTPUT: out_172 
* OUTPUT: out_173 
* OUTPUT: out_174 
* OUTPUT: out_175 
* OUTPUT: out_176 
* OUTPUT: out_177 
* OUTPUT: out_178 
* OUTPUT: out_179 
* OUTPUT: out_180 
* OUTPUT: out_181 
* OUTPUT: out_182 
* OUTPUT: out_183 
* POWER : vdd 
* GROUND: gnd 
* rows: 184 Buffer size of: 4
Xwld0
+ in_0 out_0 vdd gnd
+ sram_pinv_dec_3
Xwld1
+ in_1 out_1 vdd gnd
+ sram_pinv_dec_3
Xwld2
+ in_2 out_2 vdd gnd
+ sram_pinv_dec_3
Xwld3
+ in_3 out_3 vdd gnd
+ sram_pinv_dec_3
Xwld4
+ in_4 out_4 vdd gnd
+ sram_pinv_dec_3
Xwld5
+ in_5 out_5 vdd gnd
+ sram_pinv_dec_3
Xwld6
+ in_6 out_6 vdd gnd
+ sram_pinv_dec_3
Xwld7
+ in_7 out_7 vdd gnd
+ sram_pinv_dec_3
Xwld8
+ in_8 out_8 vdd gnd
+ sram_pinv_dec_3
Xwld9
+ in_9 out_9 vdd gnd
+ sram_pinv_dec_3
Xwld10
+ in_10 out_10 vdd gnd
+ sram_pinv_dec_3
Xwld11
+ in_11 out_11 vdd gnd
+ sram_pinv_dec_3
Xwld12
+ in_12 out_12 vdd gnd
+ sram_pinv_dec_3
Xwld13
+ in_13 out_13 vdd gnd
+ sram_pinv_dec_3
Xwld14
+ in_14 out_14 vdd gnd
+ sram_pinv_dec_3
Xwld15
+ in_15 out_15 vdd gnd
+ sram_pinv_dec_3
Xwld16
+ in_16 out_16 vdd gnd
+ sram_pinv_dec_3
Xwld17
+ in_17 out_17 vdd gnd
+ sram_pinv_dec_3
Xwld18
+ in_18 out_18 vdd gnd
+ sram_pinv_dec_3
Xwld19
+ in_19 out_19 vdd gnd
+ sram_pinv_dec_3
Xwld20
+ in_20 out_20 vdd gnd
+ sram_pinv_dec_3
Xwld21
+ in_21 out_21 vdd gnd
+ sram_pinv_dec_3
Xwld22
+ in_22 out_22 vdd gnd
+ sram_pinv_dec_3
Xwld23
+ in_23 out_23 vdd gnd
+ sram_pinv_dec_3
Xwld24
+ in_24 out_24 vdd gnd
+ sram_pinv_dec_3
Xwld25
+ in_25 out_25 vdd gnd
+ sram_pinv_dec_3
Xwld26
+ in_26 out_26 vdd gnd
+ sram_pinv_dec_3
Xwld27
+ in_27 out_27 vdd gnd
+ sram_pinv_dec_3
Xwld28
+ in_28 out_28 vdd gnd
+ sram_pinv_dec_3
Xwld29
+ in_29 out_29 vdd gnd
+ sram_pinv_dec_3
Xwld30
+ in_30 out_30 vdd gnd
+ sram_pinv_dec_3
Xwld31
+ in_31 out_31 vdd gnd
+ sram_pinv_dec_3
Xwld32
+ in_32 out_32 vdd gnd
+ sram_pinv_dec_3
Xwld33
+ in_33 out_33 vdd gnd
+ sram_pinv_dec_3
Xwld34
+ in_34 out_34 vdd gnd
+ sram_pinv_dec_3
Xwld35
+ in_35 out_35 vdd gnd
+ sram_pinv_dec_3
Xwld36
+ in_36 out_36 vdd gnd
+ sram_pinv_dec_3
Xwld37
+ in_37 out_37 vdd gnd
+ sram_pinv_dec_3
Xwld38
+ in_38 out_38 vdd gnd
+ sram_pinv_dec_3
Xwld39
+ in_39 out_39 vdd gnd
+ sram_pinv_dec_3
Xwld40
+ in_40 out_40 vdd gnd
+ sram_pinv_dec_3
Xwld41
+ in_41 out_41 vdd gnd
+ sram_pinv_dec_3
Xwld42
+ in_42 out_42 vdd gnd
+ sram_pinv_dec_3
Xwld43
+ in_43 out_43 vdd gnd
+ sram_pinv_dec_3
Xwld44
+ in_44 out_44 vdd gnd
+ sram_pinv_dec_3
Xwld45
+ in_45 out_45 vdd gnd
+ sram_pinv_dec_3
Xwld46
+ in_46 out_46 vdd gnd
+ sram_pinv_dec_3
Xwld47
+ in_47 out_47 vdd gnd
+ sram_pinv_dec_3
Xwld48
+ in_48 out_48 vdd gnd
+ sram_pinv_dec_3
Xwld49
+ in_49 out_49 vdd gnd
+ sram_pinv_dec_3
Xwld50
+ in_50 out_50 vdd gnd
+ sram_pinv_dec_3
Xwld51
+ in_51 out_51 vdd gnd
+ sram_pinv_dec_3
Xwld52
+ in_52 out_52 vdd gnd
+ sram_pinv_dec_3
Xwld53
+ in_53 out_53 vdd gnd
+ sram_pinv_dec_3
Xwld54
+ in_54 out_54 vdd gnd
+ sram_pinv_dec_3
Xwld55
+ in_55 out_55 vdd gnd
+ sram_pinv_dec_3
Xwld56
+ in_56 out_56 vdd gnd
+ sram_pinv_dec_3
Xwld57
+ in_57 out_57 vdd gnd
+ sram_pinv_dec_3
Xwld58
+ in_58 out_58 vdd gnd
+ sram_pinv_dec_3
Xwld59
+ in_59 out_59 vdd gnd
+ sram_pinv_dec_3
Xwld60
+ in_60 out_60 vdd gnd
+ sram_pinv_dec_3
Xwld61
+ in_61 out_61 vdd gnd
+ sram_pinv_dec_3
Xwld62
+ in_62 out_62 vdd gnd
+ sram_pinv_dec_3
Xwld63
+ in_63 out_63 vdd gnd
+ sram_pinv_dec_3
Xwld64
+ in_64 out_64 vdd gnd
+ sram_pinv_dec_3
Xwld65
+ in_65 out_65 vdd gnd
+ sram_pinv_dec_3
Xwld66
+ in_66 out_66 vdd gnd
+ sram_pinv_dec_3
Xwld67
+ in_67 out_67 vdd gnd
+ sram_pinv_dec_3
Xwld68
+ in_68 out_68 vdd gnd
+ sram_pinv_dec_3
Xwld69
+ in_69 out_69 vdd gnd
+ sram_pinv_dec_3
Xwld70
+ in_70 out_70 vdd gnd
+ sram_pinv_dec_3
Xwld71
+ in_71 out_71 vdd gnd
+ sram_pinv_dec_3
Xwld72
+ in_72 out_72 vdd gnd
+ sram_pinv_dec_3
Xwld73
+ in_73 out_73 vdd gnd
+ sram_pinv_dec_3
Xwld74
+ in_74 out_74 vdd gnd
+ sram_pinv_dec_3
Xwld75
+ in_75 out_75 vdd gnd
+ sram_pinv_dec_3
Xwld76
+ in_76 out_76 vdd gnd
+ sram_pinv_dec_3
Xwld77
+ in_77 out_77 vdd gnd
+ sram_pinv_dec_3
Xwld78
+ in_78 out_78 vdd gnd
+ sram_pinv_dec_3
Xwld79
+ in_79 out_79 vdd gnd
+ sram_pinv_dec_3
Xwld80
+ in_80 out_80 vdd gnd
+ sram_pinv_dec_3
Xwld81
+ in_81 out_81 vdd gnd
+ sram_pinv_dec_3
Xwld82
+ in_82 out_82 vdd gnd
+ sram_pinv_dec_3
Xwld83
+ in_83 out_83 vdd gnd
+ sram_pinv_dec_3
Xwld84
+ in_84 out_84 vdd gnd
+ sram_pinv_dec_3
Xwld85
+ in_85 out_85 vdd gnd
+ sram_pinv_dec_3
Xwld86
+ in_86 out_86 vdd gnd
+ sram_pinv_dec_3
Xwld87
+ in_87 out_87 vdd gnd
+ sram_pinv_dec_3
Xwld88
+ in_88 out_88 vdd gnd
+ sram_pinv_dec_3
Xwld89
+ in_89 out_89 vdd gnd
+ sram_pinv_dec_3
Xwld90
+ in_90 out_90 vdd gnd
+ sram_pinv_dec_3
Xwld91
+ in_91 out_91 vdd gnd
+ sram_pinv_dec_3
Xwld92
+ in_92 out_92 vdd gnd
+ sram_pinv_dec_3
Xwld93
+ in_93 out_93 vdd gnd
+ sram_pinv_dec_3
Xwld94
+ in_94 out_94 vdd gnd
+ sram_pinv_dec_3
Xwld95
+ in_95 out_95 vdd gnd
+ sram_pinv_dec_3
Xwld96
+ in_96 out_96 vdd gnd
+ sram_pinv_dec_3
Xwld97
+ in_97 out_97 vdd gnd
+ sram_pinv_dec_3
Xwld98
+ in_98 out_98 vdd gnd
+ sram_pinv_dec_3
Xwld99
+ in_99 out_99 vdd gnd
+ sram_pinv_dec_3
Xwld100
+ in_100 out_100 vdd gnd
+ sram_pinv_dec_3
Xwld101
+ in_101 out_101 vdd gnd
+ sram_pinv_dec_3
Xwld102
+ in_102 out_102 vdd gnd
+ sram_pinv_dec_3
Xwld103
+ in_103 out_103 vdd gnd
+ sram_pinv_dec_3
Xwld104
+ in_104 out_104 vdd gnd
+ sram_pinv_dec_3
Xwld105
+ in_105 out_105 vdd gnd
+ sram_pinv_dec_3
Xwld106
+ in_106 out_106 vdd gnd
+ sram_pinv_dec_3
Xwld107
+ in_107 out_107 vdd gnd
+ sram_pinv_dec_3
Xwld108
+ in_108 out_108 vdd gnd
+ sram_pinv_dec_3
Xwld109
+ in_109 out_109 vdd gnd
+ sram_pinv_dec_3
Xwld110
+ in_110 out_110 vdd gnd
+ sram_pinv_dec_3
Xwld111
+ in_111 out_111 vdd gnd
+ sram_pinv_dec_3
Xwld112
+ in_112 out_112 vdd gnd
+ sram_pinv_dec_3
Xwld113
+ in_113 out_113 vdd gnd
+ sram_pinv_dec_3
Xwld114
+ in_114 out_114 vdd gnd
+ sram_pinv_dec_3
Xwld115
+ in_115 out_115 vdd gnd
+ sram_pinv_dec_3
Xwld116
+ in_116 out_116 vdd gnd
+ sram_pinv_dec_3
Xwld117
+ in_117 out_117 vdd gnd
+ sram_pinv_dec_3
Xwld118
+ in_118 out_118 vdd gnd
+ sram_pinv_dec_3
Xwld119
+ in_119 out_119 vdd gnd
+ sram_pinv_dec_3
Xwld120
+ in_120 out_120 vdd gnd
+ sram_pinv_dec_3
Xwld121
+ in_121 out_121 vdd gnd
+ sram_pinv_dec_3
Xwld122
+ in_122 out_122 vdd gnd
+ sram_pinv_dec_3
Xwld123
+ in_123 out_123 vdd gnd
+ sram_pinv_dec_3
Xwld124
+ in_124 out_124 vdd gnd
+ sram_pinv_dec_3
Xwld125
+ in_125 out_125 vdd gnd
+ sram_pinv_dec_3
Xwld126
+ in_126 out_126 vdd gnd
+ sram_pinv_dec_3
Xwld127
+ in_127 out_127 vdd gnd
+ sram_pinv_dec_3
Xwld128
+ in_128 out_128 vdd gnd
+ sram_pinv_dec_3
Xwld129
+ in_129 out_129 vdd gnd
+ sram_pinv_dec_3
Xwld130
+ in_130 out_130 vdd gnd
+ sram_pinv_dec_3
Xwld131
+ in_131 out_131 vdd gnd
+ sram_pinv_dec_3
Xwld132
+ in_132 out_132 vdd gnd
+ sram_pinv_dec_3
Xwld133
+ in_133 out_133 vdd gnd
+ sram_pinv_dec_3
Xwld134
+ in_134 out_134 vdd gnd
+ sram_pinv_dec_3
Xwld135
+ in_135 out_135 vdd gnd
+ sram_pinv_dec_3
Xwld136
+ in_136 out_136 vdd gnd
+ sram_pinv_dec_3
Xwld137
+ in_137 out_137 vdd gnd
+ sram_pinv_dec_3
Xwld138
+ in_138 out_138 vdd gnd
+ sram_pinv_dec_3
Xwld139
+ in_139 out_139 vdd gnd
+ sram_pinv_dec_3
Xwld140
+ in_140 out_140 vdd gnd
+ sram_pinv_dec_3
Xwld141
+ in_141 out_141 vdd gnd
+ sram_pinv_dec_3
Xwld142
+ in_142 out_142 vdd gnd
+ sram_pinv_dec_3
Xwld143
+ in_143 out_143 vdd gnd
+ sram_pinv_dec_3
Xwld144
+ in_144 out_144 vdd gnd
+ sram_pinv_dec_3
Xwld145
+ in_145 out_145 vdd gnd
+ sram_pinv_dec_3
Xwld146
+ in_146 out_146 vdd gnd
+ sram_pinv_dec_3
Xwld147
+ in_147 out_147 vdd gnd
+ sram_pinv_dec_3
Xwld148
+ in_148 out_148 vdd gnd
+ sram_pinv_dec_3
Xwld149
+ in_149 out_149 vdd gnd
+ sram_pinv_dec_3
Xwld150
+ in_150 out_150 vdd gnd
+ sram_pinv_dec_3
Xwld151
+ in_151 out_151 vdd gnd
+ sram_pinv_dec_3
Xwld152
+ in_152 out_152 vdd gnd
+ sram_pinv_dec_3
Xwld153
+ in_153 out_153 vdd gnd
+ sram_pinv_dec_3
Xwld154
+ in_154 out_154 vdd gnd
+ sram_pinv_dec_3
Xwld155
+ in_155 out_155 vdd gnd
+ sram_pinv_dec_3
Xwld156
+ in_156 out_156 vdd gnd
+ sram_pinv_dec_3
Xwld157
+ in_157 out_157 vdd gnd
+ sram_pinv_dec_3
Xwld158
+ in_158 out_158 vdd gnd
+ sram_pinv_dec_3
Xwld159
+ in_159 out_159 vdd gnd
+ sram_pinv_dec_3
Xwld160
+ in_160 out_160 vdd gnd
+ sram_pinv_dec_3
Xwld161
+ in_161 out_161 vdd gnd
+ sram_pinv_dec_3
Xwld162
+ in_162 out_162 vdd gnd
+ sram_pinv_dec_3
Xwld163
+ in_163 out_163 vdd gnd
+ sram_pinv_dec_3
Xwld164
+ in_164 out_164 vdd gnd
+ sram_pinv_dec_3
Xwld165
+ in_165 out_165 vdd gnd
+ sram_pinv_dec_3
Xwld166
+ in_166 out_166 vdd gnd
+ sram_pinv_dec_3
Xwld167
+ in_167 out_167 vdd gnd
+ sram_pinv_dec_3
Xwld168
+ in_168 out_168 vdd gnd
+ sram_pinv_dec_3
Xwld169
+ in_169 out_169 vdd gnd
+ sram_pinv_dec_3
Xwld170
+ in_170 out_170 vdd gnd
+ sram_pinv_dec_3
Xwld171
+ in_171 out_171 vdd gnd
+ sram_pinv_dec_3
Xwld172
+ in_172 out_172 vdd gnd
+ sram_pinv_dec_3
Xwld173
+ in_173 out_173 vdd gnd
+ sram_pinv_dec_3
Xwld174
+ in_174 out_174 vdd gnd
+ sram_pinv_dec_3
Xwld175
+ in_175 out_175 vdd gnd
+ sram_pinv_dec_3
Xwld176
+ in_176 out_176 vdd gnd
+ sram_pinv_dec_3
Xwld177
+ in_177 out_177 vdd gnd
+ sram_pinv_dec_3
Xwld178
+ in_178 out_178 vdd gnd
+ sram_pinv_dec_3
Xwld179
+ in_179 out_179 vdd gnd
+ sram_pinv_dec_3
Xwld180
+ in_180 out_180 vdd gnd
+ sram_pinv_dec_3
Xwld181
+ in_181 out_181 vdd gnd
+ sram_pinv_dec_3
Xwld182
+ in_182 out_182 vdd gnd
+ sram_pinv_dec_3
Xwld183
+ in_183 out_183 vdd gnd
+ sram_pinv_dec_3
.ENDS sram_rom_bitline_inverter

.SUBCKT sram_pinv_dec_4
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=1.68 l=0.15 pd=3.66 ps=3.66 as=0.63u ad=0.63u
.ENDS sram_pinv_dec_4

.SUBCKT sram_rom_output_buffer
+ in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 out_0 out_1 out_2 out_3 out_4
+ out_5 out_6 out_7 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* POWER : vdd 
* GROUND: gnd 
* rows: 8 Buffer size of: 4
Xwld0
+ in_0 out_0 vdd gnd
+ sram_pinv_dec_4
Xwld1
+ in_1 out_1 vdd gnd
+ sram_pinv_dec_4
Xwld2
+ in_2 out_2 vdd gnd
+ sram_pinv_dec_4
Xwld3
+ in_3 out_3 vdd gnd
+ sram_pinv_dec_4
Xwld4
+ in_4 out_4 vdd gnd
+ sram_pinv_dec_4
Xwld5
+ in_5 out_5 vdd gnd
+ sram_pinv_dec_4
Xwld6
+ in_6 out_6 vdd gnd
+ sram_pinv_dec_4
Xwld7
+ in_7 out_7 vdd gnd
+ sram_pinv_dec_4
.ENDS sram_rom_output_buffer

.SUBCKT sram_rom_precharge_array_0
+ pre_bl0_out pre_bl1_out pre_bl2_out pre_bl3_out pre_bl4_out
+ pre_bl5_out pre_bl6_out pre_bl7_out pre_bl8_out pre_bl9_out
+ pre_bl10_out pre_bl11_out pre_bl12_out pre_bl13_out pre_bl14_out
+ pre_bl15_out pre_bl16_out pre_bl17_out pre_bl18_out pre_bl19_out
+ pre_bl20_out pre_bl21_out pre_bl22_out pre_bl23_out pre_bl24_out
+ pre_bl25_out pre_bl26_out pre_bl27_out pre_bl28_out pre_bl29_out
+ pre_bl30_out pre_bl31_out pre_bl32_out pre_bl33_out pre_bl34_out
+ pre_bl35_out pre_bl36_out pre_bl37_out pre_bl38_out pre_bl39_out
+ pre_bl40_out pre_bl41_out pre_bl42_out pre_bl43_out pre_bl44_out
+ pre_bl45_out pre_bl46_out pre_bl47_out pre_bl48_out pre_bl49_out
+ pre_bl50_out pre_bl51_out pre_bl52_out pre_bl53_out pre_bl54_out
+ pre_bl55_out pre_bl56_out pre_bl57_out pre_bl58_out pre_bl59_out
+ pre_bl60_out pre_bl61_out pre_bl62_out pre_bl63_out pre_bl64_out
+ pre_bl65_out pre_bl66_out pre_bl67_out pre_bl68_out pre_bl69_out
+ pre_bl70_out pre_bl71_out pre_bl72_out pre_bl73_out pre_bl74_out
+ pre_bl75_out pre_bl76_out pre_bl77_out pre_bl78_out pre_bl79_out
+ pre_bl80_out pre_bl81_out pre_bl82_out pre_bl83_out pre_bl84_out
+ pre_bl85_out pre_bl86_out pre_bl87_out pre_bl88_out gate vdd
* OUTPUT: pre_bl0_out 
* OUTPUT: pre_bl1_out 
* OUTPUT: pre_bl2_out 
* OUTPUT: pre_bl3_out 
* OUTPUT: pre_bl4_out 
* OUTPUT: pre_bl5_out 
* OUTPUT: pre_bl6_out 
* OUTPUT: pre_bl7_out 
* OUTPUT: pre_bl8_out 
* OUTPUT: pre_bl9_out 
* OUTPUT: pre_bl10_out 
* OUTPUT: pre_bl11_out 
* OUTPUT: pre_bl12_out 
* OUTPUT: pre_bl13_out 
* OUTPUT: pre_bl14_out 
* OUTPUT: pre_bl15_out 
* OUTPUT: pre_bl16_out 
* OUTPUT: pre_bl17_out 
* OUTPUT: pre_bl18_out 
* OUTPUT: pre_bl19_out 
* OUTPUT: pre_bl20_out 
* OUTPUT: pre_bl21_out 
* OUTPUT: pre_bl22_out 
* OUTPUT: pre_bl23_out 
* OUTPUT: pre_bl24_out 
* OUTPUT: pre_bl25_out 
* OUTPUT: pre_bl26_out 
* OUTPUT: pre_bl27_out 
* OUTPUT: pre_bl28_out 
* OUTPUT: pre_bl29_out 
* OUTPUT: pre_bl30_out 
* OUTPUT: pre_bl31_out 
* OUTPUT: pre_bl32_out 
* OUTPUT: pre_bl33_out 
* OUTPUT: pre_bl34_out 
* OUTPUT: pre_bl35_out 
* OUTPUT: pre_bl36_out 
* OUTPUT: pre_bl37_out 
* OUTPUT: pre_bl38_out 
* OUTPUT: pre_bl39_out 
* OUTPUT: pre_bl40_out 
* OUTPUT: pre_bl41_out 
* OUTPUT: pre_bl42_out 
* OUTPUT: pre_bl43_out 
* OUTPUT: pre_bl44_out 
* OUTPUT: pre_bl45_out 
* OUTPUT: pre_bl46_out 
* OUTPUT: pre_bl47_out 
* OUTPUT: pre_bl48_out 
* OUTPUT: pre_bl49_out 
* OUTPUT: pre_bl50_out 
* OUTPUT: pre_bl51_out 
* OUTPUT: pre_bl52_out 
* OUTPUT: pre_bl53_out 
* OUTPUT: pre_bl54_out 
* OUTPUT: pre_bl55_out 
* OUTPUT: pre_bl56_out 
* OUTPUT: pre_bl57_out 
* OUTPUT: pre_bl58_out 
* OUTPUT: pre_bl59_out 
* OUTPUT: pre_bl60_out 
* OUTPUT: pre_bl61_out 
* OUTPUT: pre_bl62_out 
* OUTPUT: pre_bl63_out 
* OUTPUT: pre_bl64_out 
* OUTPUT: pre_bl65_out 
* OUTPUT: pre_bl66_out 
* OUTPUT: pre_bl67_out 
* OUTPUT: pre_bl68_out 
* OUTPUT: pre_bl69_out 
* OUTPUT: pre_bl70_out 
* OUTPUT: pre_bl71_out 
* OUTPUT: pre_bl72_out 
* OUTPUT: pre_bl73_out 
* OUTPUT: pre_bl74_out 
* OUTPUT: pre_bl75_out 
* OUTPUT: pre_bl76_out 
* OUTPUT: pre_bl77_out 
* OUTPUT: pre_bl78_out 
* OUTPUT: pre_bl79_out 
* OUTPUT: pre_bl80_out 
* OUTPUT: pre_bl81_out 
* OUTPUT: pre_bl82_out 
* OUTPUT: pre_bl83_out 
* OUTPUT: pre_bl84_out 
* OUTPUT: pre_bl85_out 
* OUTPUT: pre_bl86_out 
* OUTPUT: pre_bl87_out 
* OUTPUT: pre_bl88_out 
* INPUT : gate 
* POWER : vdd 
Xpmos_c0
+ vdd gate pre_bl0_out
+ sram_precharge_cell
Xpmos_c1
+ vdd gate pre_bl1_out
+ sram_precharge_cell
Xpmos_c2
+ vdd gate pre_bl2_out
+ sram_precharge_cell
Xpmos_c3
+ vdd gate pre_bl3_out
+ sram_precharge_cell
Xpmos_c4
+ vdd gate pre_bl4_out
+ sram_precharge_cell
Xpmos_c5
+ vdd gate pre_bl5_out
+ sram_precharge_cell
Xpmos_c6
+ vdd gate pre_bl6_out
+ sram_precharge_cell
Xpmos_c7
+ vdd gate pre_bl7_out
+ sram_precharge_cell
Xpmos_c8
+ vdd gate pre_bl8_out
+ sram_precharge_cell
Xpmos_c9
+ vdd gate pre_bl9_out
+ sram_precharge_cell
Xpmos_c10
+ vdd gate pre_bl10_out
+ sram_precharge_cell
Xpmos_c11
+ vdd gate pre_bl11_out
+ sram_precharge_cell
Xpmos_c12
+ vdd gate pre_bl12_out
+ sram_precharge_cell
Xpmos_c13
+ vdd gate pre_bl13_out
+ sram_precharge_cell
Xpmos_c14
+ vdd gate pre_bl14_out
+ sram_precharge_cell
Xpmos_c15
+ vdd gate pre_bl15_out
+ sram_precharge_cell
Xpmos_c16
+ vdd gate pre_bl16_out
+ sram_precharge_cell
Xpmos_c17
+ vdd gate pre_bl17_out
+ sram_precharge_cell
Xpmos_c18
+ vdd gate pre_bl18_out
+ sram_precharge_cell
Xpmos_c19
+ vdd gate pre_bl19_out
+ sram_precharge_cell
Xpmos_c20
+ vdd gate pre_bl20_out
+ sram_precharge_cell
Xpmos_c21
+ vdd gate pre_bl21_out
+ sram_precharge_cell
Xpmos_c22
+ vdd gate pre_bl22_out
+ sram_precharge_cell
Xpmos_c23
+ vdd gate pre_bl23_out
+ sram_precharge_cell
Xpmos_c24
+ vdd gate pre_bl24_out
+ sram_precharge_cell
Xpmos_c25
+ vdd gate pre_bl25_out
+ sram_precharge_cell
Xpmos_c26
+ vdd gate pre_bl26_out
+ sram_precharge_cell
Xpmos_c27
+ vdd gate pre_bl27_out
+ sram_precharge_cell
Xpmos_c28
+ vdd gate pre_bl28_out
+ sram_precharge_cell
Xpmos_c29
+ vdd gate pre_bl29_out
+ sram_precharge_cell
Xpmos_c30
+ vdd gate pre_bl30_out
+ sram_precharge_cell
Xpmos_c31
+ vdd gate pre_bl31_out
+ sram_precharge_cell
Xpmos_c32
+ vdd gate pre_bl32_out
+ sram_precharge_cell
Xpmos_c33
+ vdd gate pre_bl33_out
+ sram_precharge_cell
Xpmos_c34
+ vdd gate pre_bl34_out
+ sram_precharge_cell
Xpmos_c35
+ vdd gate pre_bl35_out
+ sram_precharge_cell
Xpmos_c36
+ vdd gate pre_bl36_out
+ sram_precharge_cell
Xpmos_c37
+ vdd gate pre_bl37_out
+ sram_precharge_cell
Xpmos_c38
+ vdd gate pre_bl38_out
+ sram_precharge_cell
Xpmos_c39
+ vdd gate pre_bl39_out
+ sram_precharge_cell
Xpmos_c40
+ vdd gate pre_bl40_out
+ sram_precharge_cell
Xpmos_c41
+ vdd gate pre_bl41_out
+ sram_precharge_cell
Xpmos_c42
+ vdd gate pre_bl42_out
+ sram_precharge_cell
Xpmos_c43
+ vdd gate pre_bl43_out
+ sram_precharge_cell
Xpmos_c44
+ vdd gate pre_bl44_out
+ sram_precharge_cell
Xpmos_c45
+ vdd gate pre_bl45_out
+ sram_precharge_cell
Xpmos_c46
+ vdd gate pre_bl46_out
+ sram_precharge_cell
Xpmos_c47
+ vdd gate pre_bl47_out
+ sram_precharge_cell
Xpmos_c48
+ vdd gate pre_bl48_out
+ sram_precharge_cell
Xpmos_c49
+ vdd gate pre_bl49_out
+ sram_precharge_cell
Xpmos_c50
+ vdd gate pre_bl50_out
+ sram_precharge_cell
Xpmos_c51
+ vdd gate pre_bl51_out
+ sram_precharge_cell
Xpmos_c52
+ vdd gate pre_bl52_out
+ sram_precharge_cell
Xpmos_c53
+ vdd gate pre_bl53_out
+ sram_precharge_cell
Xpmos_c54
+ vdd gate pre_bl54_out
+ sram_precharge_cell
Xpmos_c55
+ vdd gate pre_bl55_out
+ sram_precharge_cell
Xpmos_c56
+ vdd gate pre_bl56_out
+ sram_precharge_cell
Xpmos_c57
+ vdd gate pre_bl57_out
+ sram_precharge_cell
Xpmos_c58
+ vdd gate pre_bl58_out
+ sram_precharge_cell
Xpmos_c59
+ vdd gate pre_bl59_out
+ sram_precharge_cell
Xpmos_c60
+ vdd gate pre_bl60_out
+ sram_precharge_cell
Xpmos_c61
+ vdd gate pre_bl61_out
+ sram_precharge_cell
Xpmos_c62
+ vdd gate pre_bl62_out
+ sram_precharge_cell
Xpmos_c63
+ vdd gate pre_bl63_out
+ sram_precharge_cell
Xpmos_c64
+ vdd gate pre_bl64_out
+ sram_precharge_cell
Xpmos_c65
+ vdd gate pre_bl65_out
+ sram_precharge_cell
Xpmos_c66
+ vdd gate pre_bl66_out
+ sram_precharge_cell
Xpmos_c67
+ vdd gate pre_bl67_out
+ sram_precharge_cell
Xpmos_c68
+ vdd gate pre_bl68_out
+ sram_precharge_cell
Xpmos_c69
+ vdd gate pre_bl69_out
+ sram_precharge_cell
Xpmos_c70
+ vdd gate pre_bl70_out
+ sram_precharge_cell
Xpmos_c71
+ vdd gate pre_bl71_out
+ sram_precharge_cell
Xpmos_c72
+ vdd gate pre_bl72_out
+ sram_precharge_cell
Xpmos_c73
+ vdd gate pre_bl73_out
+ sram_precharge_cell
Xpmos_c74
+ vdd gate pre_bl74_out
+ sram_precharge_cell
Xpmos_c75
+ vdd gate pre_bl75_out
+ sram_precharge_cell
Xpmos_c76
+ vdd gate pre_bl76_out
+ sram_precharge_cell
Xpmos_c77
+ vdd gate pre_bl77_out
+ sram_precharge_cell
Xpmos_c78
+ vdd gate pre_bl78_out
+ sram_precharge_cell
Xpmos_c79
+ vdd gate pre_bl79_out
+ sram_precharge_cell
Xpmos_c80
+ vdd gate pre_bl80_out
+ sram_precharge_cell
Xpmos_c81
+ vdd gate pre_bl81_out
+ sram_precharge_cell
Xpmos_c82
+ vdd gate pre_bl82_out
+ sram_precharge_cell
Xpmos_c83
+ vdd gate pre_bl83_out
+ sram_precharge_cell
Xpmos_c84
+ vdd gate pre_bl84_out
+ sram_precharge_cell
Xpmos_c85
+ vdd gate pre_bl85_out
+ sram_precharge_cell
Xpmos_c86
+ vdd gate pre_bl86_out
+ sram_precharge_cell
Xpmos_c87
+ vdd gate pre_bl87_out
+ sram_precharge_cell
Xpmos_c88
+ vdd gate pre_bl88_out
+ sram_precharge_cell
.ENDS sram_rom_precharge_array_0

.SUBCKT sram_rom_row_decode_array
+ bl_0_0 bl_0_1 bl_0_2 bl_0_3 bl_0_4 bl_0_5 bl_0_6 bl_0_7 bl_0_8 bl_0_9
+ bl_0_10 bl_0_11 bl_0_12 bl_0_13 bl_0_14 bl_0_15 bl_0_16 bl_0_17
+ bl_0_18 bl_0_19 bl_0_20 bl_0_21 bl_0_22 bl_0_23 bl_0_24 bl_0_25
+ bl_0_26 bl_0_27 bl_0_28 bl_0_29 bl_0_30 bl_0_31 bl_0_32 bl_0_33
+ bl_0_34 bl_0_35 bl_0_36 bl_0_37 bl_0_38 bl_0_39 bl_0_40 bl_0_41
+ bl_0_42 bl_0_43 bl_0_44 bl_0_45 bl_0_46 bl_0_47 bl_0_48 bl_0_49
+ bl_0_50 bl_0_51 bl_0_52 bl_0_53 bl_0_54 bl_0_55 bl_0_56 bl_0_57
+ bl_0_58 bl_0_59 bl_0_60 bl_0_61 bl_0_62 bl_0_63 bl_0_64 bl_0_65
+ bl_0_66 bl_0_67 bl_0_68 bl_0_69 bl_0_70 bl_0_71 bl_0_72 bl_0_73
+ bl_0_74 bl_0_75 bl_0_76 bl_0_77 bl_0_78 bl_0_79 bl_0_80 bl_0_81
+ bl_0_82 bl_0_83 bl_0_84 bl_0_85 bl_0_86 bl_0_87 bl_0_88 wl_0_0 wl_0_1
+ wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7 wl_0_8 wl_0_9 wl_0_10
+ wl_0_11 wl_0_12 wl_0_13 precharge vdd gnd
* OUTPUT: bl_0_0 
* OUTPUT: bl_0_1 
* OUTPUT: bl_0_2 
* OUTPUT: bl_0_3 
* OUTPUT: bl_0_4 
* OUTPUT: bl_0_5 
* OUTPUT: bl_0_6 
* OUTPUT: bl_0_7 
* OUTPUT: bl_0_8 
* OUTPUT: bl_0_9 
* OUTPUT: bl_0_10 
* OUTPUT: bl_0_11 
* OUTPUT: bl_0_12 
* OUTPUT: bl_0_13 
* OUTPUT: bl_0_14 
* OUTPUT: bl_0_15 
* OUTPUT: bl_0_16 
* OUTPUT: bl_0_17 
* OUTPUT: bl_0_18 
* OUTPUT: bl_0_19 
* OUTPUT: bl_0_20 
* OUTPUT: bl_0_21 
* OUTPUT: bl_0_22 
* OUTPUT: bl_0_23 
* OUTPUT: bl_0_24 
* OUTPUT: bl_0_25 
* OUTPUT: bl_0_26 
* OUTPUT: bl_0_27 
* OUTPUT: bl_0_28 
* OUTPUT: bl_0_29 
* OUTPUT: bl_0_30 
* OUTPUT: bl_0_31 
* OUTPUT: bl_0_32 
* OUTPUT: bl_0_33 
* OUTPUT: bl_0_34 
* OUTPUT: bl_0_35 
* OUTPUT: bl_0_36 
* OUTPUT: bl_0_37 
* OUTPUT: bl_0_38 
* OUTPUT: bl_0_39 
* OUTPUT: bl_0_40 
* OUTPUT: bl_0_41 
* OUTPUT: bl_0_42 
* OUTPUT: bl_0_43 
* OUTPUT: bl_0_44 
* OUTPUT: bl_0_45 
* OUTPUT: bl_0_46 
* OUTPUT: bl_0_47 
* OUTPUT: bl_0_48 
* OUTPUT: bl_0_49 
* OUTPUT: bl_0_50 
* OUTPUT: bl_0_51 
* OUTPUT: bl_0_52 
* OUTPUT: bl_0_53 
* OUTPUT: bl_0_54 
* OUTPUT: bl_0_55 
* OUTPUT: bl_0_56 
* OUTPUT: bl_0_57 
* OUTPUT: bl_0_58 
* OUTPUT: bl_0_59 
* OUTPUT: bl_0_60 
* OUTPUT: bl_0_61 
* OUTPUT: bl_0_62 
* OUTPUT: bl_0_63 
* OUTPUT: bl_0_64 
* OUTPUT: bl_0_65 
* OUTPUT: bl_0_66 
* OUTPUT: bl_0_67 
* OUTPUT: bl_0_68 
* OUTPUT: bl_0_69 
* OUTPUT: bl_0_70 
* OUTPUT: bl_0_71 
* OUTPUT: bl_0_72 
* OUTPUT: bl_0_73 
* OUTPUT: bl_0_74 
* OUTPUT: bl_0_75 
* OUTPUT: bl_0_76 
* OUTPUT: bl_0_77 
* OUTPUT: bl_0_78 
* OUTPUT: bl_0_79 
* OUTPUT: bl_0_80 
* OUTPUT: bl_0_81 
* OUTPUT: bl_0_82 
* OUTPUT: bl_0_83 
* OUTPUT: bl_0_84 
* OUTPUT: bl_0_85 
* OUTPUT: bl_0_86 
* OUTPUT: bl_0_87 
* OUTPUT: bl_0_88 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : precharge 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_int_0_0 bl_0_0 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c1
+ bl_int_0_1 bl_0_1 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c2
+ bl_int_0_2 bl_0_2 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c3
+ bl_int_0_3 bl_0_3 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c4
+ bl_int_0_4 bl_0_4 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c5
+ bl_int_0_5 bl_0_5 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c6
+ bl_int_0_6 bl_0_6 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c7
+ bl_int_0_7 bl_0_7 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c8
+ bl_int_0_8 bl_0_8 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c9
+ bl_int_0_9 bl_0_9 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c10
+ bl_int_0_10 bl_0_10 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c11
+ bl_int_0_11 bl_0_11 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c12
+ bl_int_0_12 bl_0_12 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c13
+ bl_int_0_13 bl_0_13 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c14
+ bl_int_0_14 bl_0_14 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c15
+ bl_int_0_15 bl_0_15 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c16
+ bl_int_0_16 bl_0_16 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c17
+ bl_int_0_17 bl_0_17 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c18
+ bl_int_0_18 bl_0_18 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c19
+ bl_int_0_19 bl_0_19 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c20
+ bl_int_0_20 bl_0_20 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c21
+ bl_int_0_21 bl_0_21 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c22
+ bl_int_0_22 bl_0_22 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c23
+ bl_int_0_23 bl_0_23 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c24
+ bl_int_0_24 bl_0_24 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c25
+ bl_int_0_25 bl_0_25 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c26
+ bl_int_0_26 bl_0_26 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c27
+ bl_int_0_27 bl_0_27 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c28
+ bl_int_0_28 bl_0_28 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c29
+ bl_int_0_29 bl_0_29 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c30
+ bl_int_0_30 bl_0_30 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c31
+ bl_int_0_31 bl_0_31 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c32
+ bl_int_0_32 bl_0_32 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c33
+ bl_int_0_33 bl_0_33 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c34
+ bl_int_0_34 bl_0_34 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c35
+ bl_int_0_35 bl_0_35 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c36
+ bl_int_0_36 bl_0_36 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c37
+ bl_int_0_37 bl_0_37 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c38
+ bl_int_0_38 bl_0_38 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c39
+ bl_int_0_39 bl_0_39 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c40
+ bl_int_0_40 bl_0_40 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c41
+ bl_int_0_41 bl_0_41 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c42
+ bl_int_0_42 bl_0_42 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c43
+ bl_int_0_43 bl_0_43 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c44
+ bl_int_0_44 bl_0_44 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c45
+ bl_int_0_45 bl_0_45 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c46
+ bl_int_0_46 bl_0_46 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c47
+ bl_int_0_47 bl_0_47 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c48
+ bl_int_0_48 bl_0_48 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c49
+ bl_int_0_49 bl_0_49 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c50
+ bl_int_0_50 bl_0_50 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c51
+ bl_int_0_51 bl_0_51 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c52
+ bl_int_0_52 bl_0_52 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c53
+ bl_int_0_53 bl_0_53 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c54
+ bl_int_0_54 bl_0_54 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c55
+ bl_int_0_55 bl_0_55 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c56
+ bl_int_0_56 bl_0_56 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c57
+ bl_int_0_57 bl_0_57 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c58
+ bl_int_0_58 bl_0_58 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c59
+ bl_int_0_59 bl_0_59 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c60
+ bl_int_0_60 bl_0_60 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c61
+ bl_int_0_61 bl_0_61 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c62
+ bl_int_0_62 bl_0_62 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c63
+ bl_int_0_63 bl_0_63 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c64
+ bl_0_64 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c65
+ bl_0_65 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c66
+ bl_0_66 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c67
+ bl_0_67 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c68
+ bl_0_68 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c69
+ bl_0_69 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c70
+ bl_0_70 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c71
+ bl_0_71 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c72
+ bl_0_72 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c73
+ bl_0_73 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c74
+ bl_0_74 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c75
+ bl_0_75 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c76
+ bl_0_76 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c77
+ bl_0_77 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c78
+ bl_0_78 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c79
+ bl_0_79 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c80
+ bl_0_80 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c81
+ bl_0_81 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c82
+ bl_0_82 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c83
+ bl_0_83 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c84
+ bl_0_84 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c85
+ bl_0_85 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c86
+ bl_0_86 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c87
+ bl_0_87 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r0_c88
+ bl_0_88 wl_0_0 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c0
+ bl_int_0_0 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c1
+ bl_int_0_1 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c2
+ bl_int_0_2 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c3
+ bl_int_0_3 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c4
+ bl_int_0_4 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c5
+ bl_int_0_5 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c6
+ bl_int_0_6 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c7
+ bl_int_0_7 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c8
+ bl_int_0_8 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c9
+ bl_int_0_9 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c10
+ bl_int_0_10 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c11
+ bl_int_0_11 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c12
+ bl_int_0_12 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c13
+ bl_int_0_13 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c14
+ bl_int_0_14 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c15
+ bl_int_0_15 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c16
+ bl_int_0_16 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c17
+ bl_int_0_17 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c18
+ bl_int_0_18 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c19
+ bl_int_0_19 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c20
+ bl_int_0_20 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c21
+ bl_int_0_21 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c22
+ bl_int_0_22 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c23
+ bl_int_0_23 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c24
+ bl_int_0_24 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c25
+ bl_int_0_25 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c26
+ bl_int_0_26 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c27
+ bl_int_0_27 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c28
+ bl_int_0_28 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c29
+ bl_int_0_29 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c30
+ bl_int_0_30 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c31
+ bl_int_0_31 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c32
+ bl_int_0_32 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c33
+ bl_int_0_33 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c34
+ bl_int_0_34 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c35
+ bl_int_0_35 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c36
+ bl_int_0_36 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c37
+ bl_int_0_37 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c38
+ bl_int_0_38 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c39
+ bl_int_0_39 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c40
+ bl_int_0_40 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c41
+ bl_int_0_41 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c42
+ bl_int_0_42 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c43
+ bl_int_0_43 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c44
+ bl_int_0_44 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c45
+ bl_int_0_45 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c46
+ bl_int_0_46 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c47
+ bl_int_0_47 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c48
+ bl_int_0_48 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c49
+ bl_int_0_49 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c50
+ bl_int_0_50 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c51
+ bl_int_0_51 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c52
+ bl_int_0_52 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c53
+ bl_int_0_53 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c54
+ bl_int_0_54 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c55
+ bl_int_0_55 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c56
+ bl_int_0_56 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c57
+ bl_int_0_57 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c58
+ bl_int_0_58 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c59
+ bl_int_0_59 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c60
+ bl_int_0_60 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c61
+ bl_int_0_61 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c62
+ bl_int_0_62 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c63
+ bl_int_0_63 wl_0_1 gnd
+ sram_rom_base_zero_cell
Xbit_r1_c64
+ bl_int_1_64 bl_0_64 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c65
+ bl_int_1_65 bl_0_65 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c66
+ bl_int_1_66 bl_0_66 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c67
+ bl_int_1_67 bl_0_67 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c68
+ bl_int_1_68 bl_0_68 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c69
+ bl_int_1_69 bl_0_69 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c70
+ bl_int_1_70 bl_0_70 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c71
+ bl_int_1_71 bl_0_71 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c72
+ bl_int_1_72 bl_0_72 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c73
+ bl_int_1_73 bl_0_73 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c74
+ bl_int_1_74 bl_0_74 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c75
+ bl_int_1_75 bl_0_75 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c76
+ bl_int_1_76 bl_0_76 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c77
+ bl_int_1_77 bl_0_77 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c78
+ bl_int_1_78 bl_0_78 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c79
+ bl_int_1_79 bl_0_79 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c80
+ bl_int_1_80 bl_0_80 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c81
+ bl_int_1_81 bl_0_81 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c82
+ bl_int_1_82 bl_0_82 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c83
+ bl_int_1_83 bl_0_83 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c84
+ bl_int_1_84 bl_0_84 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c85
+ bl_int_1_85 bl_0_85 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c86
+ bl_int_1_86 bl_0_86 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c87
+ bl_int_1_87 bl_0_87 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c88
+ bl_int_1_88 bl_0_88 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r2_c0
+ bl_int_2_0 bl_int_0_0 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c1
+ bl_int_2_1 bl_int_0_1 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c2
+ bl_int_2_2 bl_int_0_2 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c3
+ bl_int_2_3 bl_int_0_3 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c4
+ bl_int_2_4 bl_int_0_4 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c5
+ bl_int_2_5 bl_int_0_5 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c6
+ bl_int_2_6 bl_int_0_6 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c7
+ bl_int_2_7 bl_int_0_7 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c8
+ bl_int_2_8 bl_int_0_8 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c9
+ bl_int_2_9 bl_int_0_9 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c10
+ bl_int_2_10 bl_int_0_10 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c11
+ bl_int_2_11 bl_int_0_11 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c12
+ bl_int_2_12 bl_int_0_12 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c13
+ bl_int_2_13 bl_int_0_13 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c14
+ bl_int_2_14 bl_int_0_14 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c15
+ bl_int_2_15 bl_int_0_15 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c16
+ bl_int_2_16 bl_int_0_16 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c17
+ bl_int_2_17 bl_int_0_17 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c18
+ bl_int_2_18 bl_int_0_18 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c19
+ bl_int_2_19 bl_int_0_19 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c20
+ bl_int_2_20 bl_int_0_20 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c21
+ bl_int_2_21 bl_int_0_21 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c22
+ bl_int_2_22 bl_int_0_22 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c23
+ bl_int_2_23 bl_int_0_23 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c24
+ bl_int_2_24 bl_int_0_24 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c25
+ bl_int_2_25 bl_int_0_25 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c26
+ bl_int_2_26 bl_int_0_26 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c27
+ bl_int_2_27 bl_int_0_27 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c28
+ bl_int_2_28 bl_int_0_28 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c29
+ bl_int_2_29 bl_int_0_29 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c30
+ bl_int_2_30 bl_int_0_30 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c31
+ bl_int_2_31 bl_int_0_31 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c32
+ bl_int_0_32 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c33
+ bl_int_0_33 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c34
+ bl_int_0_34 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c35
+ bl_int_0_35 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c36
+ bl_int_0_36 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c37
+ bl_int_0_37 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c38
+ bl_int_0_38 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c39
+ bl_int_0_39 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c40
+ bl_int_0_40 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c41
+ bl_int_0_41 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c42
+ bl_int_0_42 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c43
+ bl_int_0_43 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c44
+ bl_int_0_44 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c45
+ bl_int_0_45 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c46
+ bl_int_0_46 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c47
+ bl_int_0_47 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c48
+ bl_int_0_48 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c49
+ bl_int_0_49 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c50
+ bl_int_0_50 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c51
+ bl_int_0_51 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c52
+ bl_int_0_52 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c53
+ bl_int_0_53 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c54
+ bl_int_0_54 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c55
+ bl_int_0_55 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c56
+ bl_int_0_56 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c57
+ bl_int_0_57 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c58
+ bl_int_0_58 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c59
+ bl_int_0_59 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c60
+ bl_int_0_60 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c61
+ bl_int_0_61 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c62
+ bl_int_0_62 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c63
+ bl_int_0_63 wl_0_2 gnd
+ sram_rom_base_zero_cell
Xbit_r2_c64
+ bl_int_2_64 bl_int_1_64 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c65
+ bl_int_2_65 bl_int_1_65 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c66
+ bl_int_2_66 bl_int_1_66 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c67
+ bl_int_2_67 bl_int_1_67 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c68
+ bl_int_2_68 bl_int_1_68 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c69
+ bl_int_2_69 bl_int_1_69 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c70
+ bl_int_2_70 bl_int_1_70 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c71
+ bl_int_2_71 bl_int_1_71 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c72
+ bl_int_2_72 bl_int_1_72 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c73
+ bl_int_2_73 bl_int_1_73 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c74
+ bl_int_2_74 bl_int_1_74 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c75
+ bl_int_2_75 bl_int_1_75 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c76
+ bl_int_2_76 bl_int_1_76 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c77
+ bl_int_2_77 bl_int_1_77 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c78
+ bl_int_2_78 bl_int_1_78 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c79
+ bl_int_2_79 bl_int_1_79 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c80
+ bl_int_2_80 bl_int_1_80 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c81
+ bl_int_2_81 bl_int_1_81 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c82
+ bl_int_2_82 bl_int_1_82 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c83
+ bl_int_2_83 bl_int_1_83 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c84
+ bl_int_2_84 bl_int_1_84 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c85
+ bl_int_2_85 bl_int_1_85 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c86
+ bl_int_2_86 bl_int_1_86 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c87
+ bl_int_2_87 bl_int_1_87 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c88
+ bl_int_2_88 bl_int_1_88 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r3_c0
+ bl_int_2_0 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c1
+ bl_int_2_1 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c2
+ bl_int_2_2 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c3
+ bl_int_2_3 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c4
+ bl_int_2_4 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c5
+ bl_int_2_5 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c6
+ bl_int_2_6 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c7
+ bl_int_2_7 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c8
+ bl_int_2_8 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c9
+ bl_int_2_9 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c10
+ bl_int_2_10 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c11
+ bl_int_2_11 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c12
+ bl_int_2_12 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c13
+ bl_int_2_13 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c14
+ bl_int_2_14 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c15
+ bl_int_2_15 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c16
+ bl_int_2_16 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c17
+ bl_int_2_17 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c18
+ bl_int_2_18 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c19
+ bl_int_2_19 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c20
+ bl_int_2_20 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c21
+ bl_int_2_21 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c22
+ bl_int_2_22 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c23
+ bl_int_2_23 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c24
+ bl_int_2_24 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c25
+ bl_int_2_25 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c26
+ bl_int_2_26 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c27
+ bl_int_2_27 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c28
+ bl_int_2_28 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c29
+ bl_int_2_29 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c30
+ bl_int_2_30 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c31
+ bl_int_2_31 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c32
+ bl_int_3_32 bl_int_0_32 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c33
+ bl_int_3_33 bl_int_0_33 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c34
+ bl_int_3_34 bl_int_0_34 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c35
+ bl_int_3_35 bl_int_0_35 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c36
+ bl_int_3_36 bl_int_0_36 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c37
+ bl_int_3_37 bl_int_0_37 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c38
+ bl_int_3_38 bl_int_0_38 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c39
+ bl_int_3_39 bl_int_0_39 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c40
+ bl_int_3_40 bl_int_0_40 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c41
+ bl_int_3_41 bl_int_0_41 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c42
+ bl_int_3_42 bl_int_0_42 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c43
+ bl_int_3_43 bl_int_0_43 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c44
+ bl_int_3_44 bl_int_0_44 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c45
+ bl_int_3_45 bl_int_0_45 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c46
+ bl_int_3_46 bl_int_0_46 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c47
+ bl_int_3_47 bl_int_0_47 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c48
+ bl_int_3_48 bl_int_0_48 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c49
+ bl_int_3_49 bl_int_0_49 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c50
+ bl_int_3_50 bl_int_0_50 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c51
+ bl_int_3_51 bl_int_0_51 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c52
+ bl_int_3_52 bl_int_0_52 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c53
+ bl_int_3_53 bl_int_0_53 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c54
+ bl_int_3_54 bl_int_0_54 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c55
+ bl_int_3_55 bl_int_0_55 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c56
+ bl_int_3_56 bl_int_0_56 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c57
+ bl_int_3_57 bl_int_0_57 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c58
+ bl_int_3_58 bl_int_0_58 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c59
+ bl_int_3_59 bl_int_0_59 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c60
+ bl_int_3_60 bl_int_0_60 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c61
+ bl_int_3_61 bl_int_0_61 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c62
+ bl_int_3_62 bl_int_0_62 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c63
+ bl_int_3_63 bl_int_0_63 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c64
+ bl_int_2_64 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c65
+ bl_int_2_65 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c66
+ bl_int_2_66 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c67
+ bl_int_2_67 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c68
+ bl_int_2_68 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c69
+ bl_int_2_69 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c70
+ bl_int_2_70 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c71
+ bl_int_2_71 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c72
+ bl_int_2_72 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c73
+ bl_int_2_73 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c74
+ bl_int_2_74 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c75
+ bl_int_2_75 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c76
+ bl_int_2_76 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c77
+ bl_int_2_77 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c78
+ bl_int_2_78 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c79
+ bl_int_2_79 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c80
+ bl_int_2_80 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c81
+ bl_int_2_81 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c82
+ bl_int_2_82 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c83
+ bl_int_2_83 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c84
+ bl_int_2_84 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c85
+ bl_int_2_85 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c86
+ bl_int_2_86 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c87
+ bl_int_2_87 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r3_c88
+ bl_int_2_88 wl_0_3 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c0
+ bl_int_4_0 bl_int_2_0 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c1
+ bl_int_4_1 bl_int_2_1 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c2
+ bl_int_4_2 bl_int_2_2 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c3
+ bl_int_4_3 bl_int_2_3 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c4
+ bl_int_4_4 bl_int_2_4 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c5
+ bl_int_4_5 bl_int_2_5 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c6
+ bl_int_4_6 bl_int_2_6 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c7
+ bl_int_4_7 bl_int_2_7 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c8
+ bl_int_4_8 bl_int_2_8 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c9
+ bl_int_4_9 bl_int_2_9 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c10
+ bl_int_4_10 bl_int_2_10 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c11
+ bl_int_4_11 bl_int_2_11 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c12
+ bl_int_4_12 bl_int_2_12 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c13
+ bl_int_4_13 bl_int_2_13 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c14
+ bl_int_4_14 bl_int_2_14 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c15
+ bl_int_4_15 bl_int_2_15 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c16
+ bl_int_2_16 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c17
+ bl_int_2_17 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c18
+ bl_int_2_18 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c19
+ bl_int_2_19 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c20
+ bl_int_2_20 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c21
+ bl_int_2_21 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c22
+ bl_int_2_22 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c23
+ bl_int_2_23 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c24
+ bl_int_2_24 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c25
+ bl_int_2_25 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c26
+ bl_int_2_26 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c27
+ bl_int_2_27 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c28
+ bl_int_2_28 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c29
+ bl_int_2_29 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c30
+ bl_int_2_30 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c31
+ bl_int_2_31 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c32
+ bl_int_4_32 bl_int_3_32 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c33
+ bl_int_4_33 bl_int_3_33 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c34
+ bl_int_4_34 bl_int_3_34 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c35
+ bl_int_4_35 bl_int_3_35 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c36
+ bl_int_4_36 bl_int_3_36 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c37
+ bl_int_4_37 bl_int_3_37 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c38
+ bl_int_4_38 bl_int_3_38 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c39
+ bl_int_4_39 bl_int_3_39 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c40
+ bl_int_4_40 bl_int_3_40 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c41
+ bl_int_4_41 bl_int_3_41 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c42
+ bl_int_4_42 bl_int_3_42 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c43
+ bl_int_4_43 bl_int_3_43 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c44
+ bl_int_4_44 bl_int_3_44 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c45
+ bl_int_4_45 bl_int_3_45 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c46
+ bl_int_4_46 bl_int_3_46 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c47
+ bl_int_4_47 bl_int_3_47 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c48
+ bl_int_3_48 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c49
+ bl_int_3_49 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c50
+ bl_int_3_50 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c51
+ bl_int_3_51 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c52
+ bl_int_3_52 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c53
+ bl_int_3_53 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c54
+ bl_int_3_54 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c55
+ bl_int_3_55 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c56
+ bl_int_3_56 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c57
+ bl_int_3_57 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c58
+ bl_int_3_58 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c59
+ bl_int_3_59 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c60
+ bl_int_3_60 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c61
+ bl_int_3_61 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c62
+ bl_int_3_62 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c63
+ bl_int_3_63 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c64
+ bl_int_4_64 bl_int_2_64 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c65
+ bl_int_4_65 bl_int_2_65 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c66
+ bl_int_4_66 bl_int_2_66 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c67
+ bl_int_4_67 bl_int_2_67 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c68
+ bl_int_4_68 bl_int_2_68 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c69
+ bl_int_4_69 bl_int_2_69 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c70
+ bl_int_4_70 bl_int_2_70 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c71
+ bl_int_4_71 bl_int_2_71 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c72
+ bl_int_4_72 bl_int_2_72 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c73
+ bl_int_4_73 bl_int_2_73 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c74
+ bl_int_4_74 bl_int_2_74 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c75
+ bl_int_4_75 bl_int_2_75 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c76
+ bl_int_4_76 bl_int_2_76 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c77
+ bl_int_4_77 bl_int_2_77 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c78
+ bl_int_4_78 bl_int_2_78 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c79
+ bl_int_4_79 bl_int_2_79 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c80
+ bl_int_2_80 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c81
+ bl_int_2_81 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c82
+ bl_int_2_82 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c83
+ bl_int_2_83 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c84
+ bl_int_2_84 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c85
+ bl_int_2_85 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c86
+ bl_int_2_86 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c87
+ bl_int_2_87 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r4_c88
+ bl_int_2_88 wl_0_4 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c0
+ bl_int_4_0 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c1
+ bl_int_4_1 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c2
+ bl_int_4_2 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c3
+ bl_int_4_3 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c4
+ bl_int_4_4 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c5
+ bl_int_4_5 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c6
+ bl_int_4_6 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c7
+ bl_int_4_7 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c8
+ bl_int_4_8 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c9
+ bl_int_4_9 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c10
+ bl_int_4_10 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c11
+ bl_int_4_11 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c12
+ bl_int_4_12 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c13
+ bl_int_4_13 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c14
+ bl_int_4_14 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c15
+ bl_int_4_15 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c16
+ bl_int_5_16 bl_int_2_16 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c17
+ bl_int_5_17 bl_int_2_17 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c18
+ bl_int_5_18 bl_int_2_18 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c19
+ bl_int_5_19 bl_int_2_19 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c20
+ bl_int_5_20 bl_int_2_20 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c21
+ bl_int_5_21 bl_int_2_21 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c22
+ bl_int_5_22 bl_int_2_22 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c23
+ bl_int_5_23 bl_int_2_23 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c24
+ bl_int_5_24 bl_int_2_24 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c25
+ bl_int_5_25 bl_int_2_25 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c26
+ bl_int_5_26 bl_int_2_26 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c27
+ bl_int_5_27 bl_int_2_27 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c28
+ bl_int_5_28 bl_int_2_28 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c29
+ bl_int_5_29 bl_int_2_29 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c30
+ bl_int_5_30 bl_int_2_30 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c31
+ bl_int_5_31 bl_int_2_31 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c32
+ bl_int_4_32 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c33
+ bl_int_4_33 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c34
+ bl_int_4_34 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c35
+ bl_int_4_35 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c36
+ bl_int_4_36 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c37
+ bl_int_4_37 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c38
+ bl_int_4_38 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c39
+ bl_int_4_39 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c40
+ bl_int_4_40 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c41
+ bl_int_4_41 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c42
+ bl_int_4_42 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c43
+ bl_int_4_43 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c44
+ bl_int_4_44 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c45
+ bl_int_4_45 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c46
+ bl_int_4_46 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c47
+ bl_int_4_47 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c48
+ bl_int_5_48 bl_int_3_48 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c49
+ bl_int_5_49 bl_int_3_49 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c50
+ bl_int_5_50 bl_int_3_50 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c51
+ bl_int_5_51 bl_int_3_51 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c52
+ bl_int_5_52 bl_int_3_52 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c53
+ bl_int_5_53 bl_int_3_53 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c54
+ bl_int_5_54 bl_int_3_54 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c55
+ bl_int_5_55 bl_int_3_55 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c56
+ bl_int_5_56 bl_int_3_56 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c57
+ bl_int_5_57 bl_int_3_57 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c58
+ bl_int_5_58 bl_int_3_58 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c59
+ bl_int_5_59 bl_int_3_59 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c60
+ bl_int_5_60 bl_int_3_60 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c61
+ bl_int_5_61 bl_int_3_61 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c62
+ bl_int_5_62 bl_int_3_62 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c63
+ bl_int_5_63 bl_int_3_63 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c64
+ bl_int_4_64 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c65
+ bl_int_4_65 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c66
+ bl_int_4_66 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c67
+ bl_int_4_67 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c68
+ bl_int_4_68 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c69
+ bl_int_4_69 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c70
+ bl_int_4_70 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c71
+ bl_int_4_71 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c72
+ bl_int_4_72 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c73
+ bl_int_4_73 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c74
+ bl_int_4_74 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c75
+ bl_int_4_75 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c76
+ bl_int_4_76 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c77
+ bl_int_4_77 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c78
+ bl_int_4_78 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c79
+ bl_int_4_79 wl_0_5 gnd
+ sram_rom_base_zero_cell
Xbit_r5_c80
+ bl_int_5_80 bl_int_2_80 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c81
+ bl_int_5_81 bl_int_2_81 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c82
+ bl_int_5_82 bl_int_2_82 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c83
+ bl_int_5_83 bl_int_2_83 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c84
+ bl_int_5_84 bl_int_2_84 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c85
+ bl_int_5_85 bl_int_2_85 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c86
+ bl_int_5_86 bl_int_2_86 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c87
+ bl_int_5_87 bl_int_2_87 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c88
+ bl_int_5_88 bl_int_2_88 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r6_c0
+ bl_int_6_0 bl_int_4_0 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c1
+ bl_int_6_1 bl_int_4_1 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c2
+ bl_int_6_2 bl_int_4_2 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c3
+ bl_int_6_3 bl_int_4_3 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c4
+ bl_int_6_4 bl_int_4_4 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c5
+ bl_int_6_5 bl_int_4_5 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c6
+ bl_int_6_6 bl_int_4_6 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c7
+ bl_int_6_7 bl_int_4_7 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c8
+ bl_int_4_8 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c9
+ bl_int_4_9 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c10
+ bl_int_4_10 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c11
+ bl_int_4_11 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c12
+ bl_int_4_12 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c13
+ bl_int_4_13 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c14
+ bl_int_4_14 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c15
+ bl_int_4_15 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c16
+ bl_int_6_16 bl_int_5_16 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c17
+ bl_int_6_17 bl_int_5_17 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c18
+ bl_int_6_18 bl_int_5_18 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c19
+ bl_int_6_19 bl_int_5_19 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c20
+ bl_int_6_20 bl_int_5_20 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c21
+ bl_int_6_21 bl_int_5_21 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c22
+ bl_int_6_22 bl_int_5_22 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c23
+ bl_int_6_23 bl_int_5_23 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c24
+ bl_int_5_24 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c25
+ bl_int_5_25 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c26
+ bl_int_5_26 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c27
+ bl_int_5_27 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c28
+ bl_int_5_28 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c29
+ bl_int_5_29 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c30
+ bl_int_5_30 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c31
+ bl_int_5_31 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c32
+ bl_int_6_32 bl_int_4_32 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c33
+ bl_int_6_33 bl_int_4_33 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c34
+ bl_int_6_34 bl_int_4_34 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c35
+ bl_int_6_35 bl_int_4_35 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c36
+ bl_int_6_36 bl_int_4_36 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c37
+ bl_int_6_37 bl_int_4_37 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c38
+ bl_int_6_38 bl_int_4_38 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c39
+ bl_int_6_39 bl_int_4_39 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c40
+ bl_int_4_40 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c41
+ bl_int_4_41 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c42
+ bl_int_4_42 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c43
+ bl_int_4_43 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c44
+ bl_int_4_44 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c45
+ bl_int_4_45 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c46
+ bl_int_4_46 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c47
+ bl_int_4_47 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c48
+ bl_int_6_48 bl_int_5_48 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c49
+ bl_int_6_49 bl_int_5_49 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c50
+ bl_int_6_50 bl_int_5_50 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c51
+ bl_int_6_51 bl_int_5_51 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c52
+ bl_int_6_52 bl_int_5_52 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c53
+ bl_int_6_53 bl_int_5_53 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c54
+ bl_int_6_54 bl_int_5_54 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c55
+ bl_int_6_55 bl_int_5_55 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c56
+ bl_int_5_56 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c57
+ bl_int_5_57 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c58
+ bl_int_5_58 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c59
+ bl_int_5_59 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c60
+ bl_int_5_60 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c61
+ bl_int_5_61 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c62
+ bl_int_5_62 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c63
+ bl_int_5_63 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c64
+ bl_int_6_64 bl_int_4_64 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c65
+ bl_int_6_65 bl_int_4_65 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c66
+ bl_int_6_66 bl_int_4_66 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c67
+ bl_int_6_67 bl_int_4_67 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c68
+ bl_int_6_68 bl_int_4_68 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c69
+ bl_int_6_69 bl_int_4_69 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c70
+ bl_int_6_70 bl_int_4_70 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c71
+ bl_int_6_71 bl_int_4_71 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c72
+ bl_int_4_72 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c73
+ bl_int_4_73 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c74
+ bl_int_4_74 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c75
+ bl_int_4_75 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c76
+ bl_int_4_76 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c77
+ bl_int_4_77 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c78
+ bl_int_4_78 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c79
+ bl_int_4_79 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r6_c80
+ bl_int_6_80 bl_int_5_80 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c81
+ bl_int_6_81 bl_int_5_81 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c82
+ bl_int_6_82 bl_int_5_82 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c83
+ bl_int_6_83 bl_int_5_83 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c84
+ bl_int_6_84 bl_int_5_84 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c85
+ bl_int_6_85 bl_int_5_85 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c86
+ bl_int_6_86 bl_int_5_86 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c87
+ bl_int_6_87 bl_int_5_87 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c88
+ bl_int_5_88 wl_0_6 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c0
+ bl_int_6_0 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c1
+ bl_int_6_1 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c2
+ bl_int_6_2 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c3
+ bl_int_6_3 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c4
+ bl_int_6_4 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c5
+ bl_int_6_5 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c6
+ bl_int_6_6 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c7
+ bl_int_6_7 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c8
+ bl_int_7_8 bl_int_4_8 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c9
+ bl_int_7_9 bl_int_4_9 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c10
+ bl_int_7_10 bl_int_4_10 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c11
+ bl_int_7_11 bl_int_4_11 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c12
+ bl_int_7_12 bl_int_4_12 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c13
+ bl_int_7_13 bl_int_4_13 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c14
+ bl_int_7_14 bl_int_4_14 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c15
+ bl_int_7_15 bl_int_4_15 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c16
+ bl_int_6_16 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c17
+ bl_int_6_17 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c18
+ bl_int_6_18 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c19
+ bl_int_6_19 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c20
+ bl_int_6_20 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c21
+ bl_int_6_21 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c22
+ bl_int_6_22 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c23
+ bl_int_6_23 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c24
+ bl_int_7_24 bl_int_5_24 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c25
+ bl_int_7_25 bl_int_5_25 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c26
+ bl_int_7_26 bl_int_5_26 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c27
+ bl_int_7_27 bl_int_5_27 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c28
+ bl_int_7_28 bl_int_5_28 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c29
+ bl_int_7_29 bl_int_5_29 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c30
+ bl_int_7_30 bl_int_5_30 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c31
+ bl_int_7_31 bl_int_5_31 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c32
+ bl_int_6_32 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c33
+ bl_int_6_33 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c34
+ bl_int_6_34 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c35
+ bl_int_6_35 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c36
+ bl_int_6_36 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c37
+ bl_int_6_37 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c38
+ bl_int_6_38 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c39
+ bl_int_6_39 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c40
+ bl_int_7_40 bl_int_4_40 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c41
+ bl_int_7_41 bl_int_4_41 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c42
+ bl_int_7_42 bl_int_4_42 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c43
+ bl_int_7_43 bl_int_4_43 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c44
+ bl_int_7_44 bl_int_4_44 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c45
+ bl_int_7_45 bl_int_4_45 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c46
+ bl_int_7_46 bl_int_4_46 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c47
+ bl_int_7_47 bl_int_4_47 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c48
+ bl_int_6_48 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c49
+ bl_int_6_49 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c50
+ bl_int_6_50 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c51
+ bl_int_6_51 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c52
+ bl_int_6_52 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c53
+ bl_int_6_53 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c54
+ bl_int_6_54 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c55
+ bl_int_6_55 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c56
+ bl_int_7_56 bl_int_5_56 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c57
+ bl_int_7_57 bl_int_5_57 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c58
+ bl_int_7_58 bl_int_5_58 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c59
+ bl_int_7_59 bl_int_5_59 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c60
+ bl_int_7_60 bl_int_5_60 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c61
+ bl_int_7_61 bl_int_5_61 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c62
+ bl_int_7_62 bl_int_5_62 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c63
+ bl_int_7_63 bl_int_5_63 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c64
+ bl_int_6_64 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c65
+ bl_int_6_65 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c66
+ bl_int_6_66 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c67
+ bl_int_6_67 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c68
+ bl_int_6_68 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c69
+ bl_int_6_69 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c70
+ bl_int_6_70 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c71
+ bl_int_6_71 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c72
+ bl_int_7_72 bl_int_4_72 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c73
+ bl_int_7_73 bl_int_4_73 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c74
+ bl_int_7_74 bl_int_4_74 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c75
+ bl_int_7_75 bl_int_4_75 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c76
+ bl_int_7_76 bl_int_4_76 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c77
+ bl_int_7_77 bl_int_4_77 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c78
+ bl_int_7_78 bl_int_4_78 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c79
+ bl_int_7_79 bl_int_4_79 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c80
+ bl_int_6_80 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c81
+ bl_int_6_81 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c82
+ bl_int_6_82 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c83
+ bl_int_6_83 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c84
+ bl_int_6_84 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c85
+ bl_int_6_85 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c86
+ bl_int_6_86 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c87
+ bl_int_6_87 wl_0_7 gnd
+ sram_rom_base_zero_cell
Xbit_r7_c88
+ bl_int_7_88 bl_int_5_88 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r8_c0
+ bl_int_8_0 bl_int_6_0 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c1
+ bl_int_8_1 bl_int_6_1 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c2
+ bl_int_8_2 bl_int_6_2 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c3
+ bl_int_8_3 bl_int_6_3 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c4
+ bl_int_6_4 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c5
+ bl_int_6_5 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c6
+ bl_int_6_6 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c7
+ bl_int_6_7 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c8
+ bl_int_8_8 bl_int_7_8 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c9
+ bl_int_8_9 bl_int_7_9 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c10
+ bl_int_8_10 bl_int_7_10 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c11
+ bl_int_8_11 bl_int_7_11 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c12
+ bl_int_7_12 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c13
+ bl_int_7_13 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c14
+ bl_int_7_14 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c15
+ bl_int_7_15 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c16
+ bl_int_8_16 bl_int_6_16 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c17
+ bl_int_8_17 bl_int_6_17 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c18
+ bl_int_8_18 bl_int_6_18 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c19
+ bl_int_8_19 bl_int_6_19 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c20
+ bl_int_6_20 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c21
+ bl_int_6_21 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c22
+ bl_int_6_22 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c23
+ bl_int_6_23 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c24
+ bl_int_8_24 bl_int_7_24 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c25
+ bl_int_8_25 bl_int_7_25 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c26
+ bl_int_8_26 bl_int_7_26 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c27
+ bl_int_8_27 bl_int_7_27 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c28
+ bl_int_7_28 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c29
+ bl_int_7_29 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c30
+ bl_int_7_30 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c31
+ bl_int_7_31 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c32
+ bl_int_8_32 bl_int_6_32 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c33
+ bl_int_8_33 bl_int_6_33 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c34
+ bl_int_8_34 bl_int_6_34 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c35
+ bl_int_8_35 bl_int_6_35 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c36
+ bl_int_6_36 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c37
+ bl_int_6_37 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c38
+ bl_int_6_38 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c39
+ bl_int_6_39 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c40
+ bl_int_8_40 bl_int_7_40 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c41
+ bl_int_8_41 bl_int_7_41 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c42
+ bl_int_8_42 bl_int_7_42 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c43
+ bl_int_8_43 bl_int_7_43 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c44
+ bl_int_7_44 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c45
+ bl_int_7_45 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c46
+ bl_int_7_46 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c47
+ bl_int_7_47 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c48
+ bl_int_8_48 bl_int_6_48 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c49
+ bl_int_8_49 bl_int_6_49 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c50
+ bl_int_8_50 bl_int_6_50 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c51
+ bl_int_8_51 bl_int_6_51 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c52
+ bl_int_6_52 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c53
+ bl_int_6_53 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c54
+ bl_int_6_54 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c55
+ bl_int_6_55 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c56
+ bl_int_8_56 bl_int_7_56 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c57
+ bl_int_8_57 bl_int_7_57 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c58
+ bl_int_8_58 bl_int_7_58 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c59
+ bl_int_8_59 bl_int_7_59 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c60
+ bl_int_7_60 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c61
+ bl_int_7_61 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c62
+ bl_int_7_62 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c63
+ bl_int_7_63 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c64
+ bl_int_8_64 bl_int_6_64 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c65
+ bl_int_8_65 bl_int_6_65 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c66
+ bl_int_8_66 bl_int_6_66 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c67
+ bl_int_8_67 bl_int_6_67 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c68
+ bl_int_6_68 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c69
+ bl_int_6_69 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c70
+ bl_int_6_70 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c71
+ bl_int_6_71 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c72
+ bl_int_8_72 bl_int_7_72 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c73
+ bl_int_8_73 bl_int_7_73 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c74
+ bl_int_8_74 bl_int_7_74 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c75
+ bl_int_8_75 bl_int_7_75 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c76
+ bl_int_7_76 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c77
+ bl_int_7_77 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c78
+ bl_int_7_78 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c79
+ bl_int_7_79 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c80
+ bl_int_8_80 bl_int_6_80 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c81
+ bl_int_8_81 bl_int_6_81 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c82
+ bl_int_8_82 bl_int_6_82 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c83
+ bl_int_8_83 bl_int_6_83 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c84
+ bl_int_6_84 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c85
+ bl_int_6_85 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c86
+ bl_int_6_86 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c87
+ bl_int_6_87 wl_0_8 gnd
+ sram_rom_base_zero_cell
Xbit_r8_c88
+ bl_int_8_88 bl_int_7_88 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r9_c0
+ bl_int_8_0 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c1
+ bl_int_8_1 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c2
+ bl_int_8_2 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c3
+ bl_int_8_3 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c4
+ bl_int_9_4 bl_int_6_4 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c5
+ bl_int_9_5 bl_int_6_5 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c6
+ bl_int_9_6 bl_int_6_6 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c7
+ bl_int_9_7 bl_int_6_7 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c8
+ bl_int_8_8 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c9
+ bl_int_8_9 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c10
+ bl_int_8_10 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c11
+ bl_int_8_11 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c12
+ bl_int_9_12 bl_int_7_12 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c13
+ bl_int_9_13 bl_int_7_13 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c14
+ bl_int_9_14 bl_int_7_14 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c15
+ bl_int_9_15 bl_int_7_15 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c16
+ bl_int_8_16 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c17
+ bl_int_8_17 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c18
+ bl_int_8_18 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c19
+ bl_int_8_19 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c20
+ bl_int_9_20 bl_int_6_20 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c21
+ bl_int_9_21 bl_int_6_21 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c22
+ bl_int_9_22 bl_int_6_22 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c23
+ bl_int_9_23 bl_int_6_23 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c24
+ bl_int_8_24 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c25
+ bl_int_8_25 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c26
+ bl_int_8_26 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c27
+ bl_int_8_27 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c28
+ bl_int_9_28 bl_int_7_28 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c29
+ bl_int_9_29 bl_int_7_29 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c30
+ bl_int_9_30 bl_int_7_30 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c31
+ bl_int_9_31 bl_int_7_31 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c32
+ bl_int_8_32 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c33
+ bl_int_8_33 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c34
+ bl_int_8_34 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c35
+ bl_int_8_35 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c36
+ bl_int_9_36 bl_int_6_36 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c37
+ bl_int_9_37 bl_int_6_37 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c38
+ bl_int_9_38 bl_int_6_38 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c39
+ bl_int_9_39 bl_int_6_39 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c40
+ bl_int_8_40 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c41
+ bl_int_8_41 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c42
+ bl_int_8_42 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c43
+ bl_int_8_43 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c44
+ bl_int_9_44 bl_int_7_44 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c45
+ bl_int_9_45 bl_int_7_45 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c46
+ bl_int_9_46 bl_int_7_46 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c47
+ bl_int_9_47 bl_int_7_47 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c48
+ bl_int_8_48 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c49
+ bl_int_8_49 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c50
+ bl_int_8_50 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c51
+ bl_int_8_51 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c52
+ bl_int_9_52 bl_int_6_52 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c53
+ bl_int_9_53 bl_int_6_53 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c54
+ bl_int_9_54 bl_int_6_54 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c55
+ bl_int_9_55 bl_int_6_55 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c56
+ bl_int_8_56 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c57
+ bl_int_8_57 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c58
+ bl_int_8_58 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c59
+ bl_int_8_59 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c60
+ bl_int_9_60 bl_int_7_60 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c61
+ bl_int_9_61 bl_int_7_61 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c62
+ bl_int_9_62 bl_int_7_62 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c63
+ bl_int_9_63 bl_int_7_63 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c64
+ bl_int_8_64 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c65
+ bl_int_8_65 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c66
+ bl_int_8_66 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c67
+ bl_int_8_67 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c68
+ bl_int_9_68 bl_int_6_68 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c69
+ bl_int_9_69 bl_int_6_69 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c70
+ bl_int_9_70 bl_int_6_70 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c71
+ bl_int_9_71 bl_int_6_71 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c72
+ bl_int_8_72 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c73
+ bl_int_8_73 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c74
+ bl_int_8_74 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c75
+ bl_int_8_75 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c76
+ bl_int_9_76 bl_int_7_76 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c77
+ bl_int_9_77 bl_int_7_77 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c78
+ bl_int_9_78 bl_int_7_78 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c79
+ bl_int_9_79 bl_int_7_79 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c80
+ bl_int_8_80 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c81
+ bl_int_8_81 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c82
+ bl_int_8_82 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c83
+ bl_int_8_83 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r9_c84
+ bl_int_9_84 bl_int_6_84 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c85
+ bl_int_9_85 bl_int_6_85 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c86
+ bl_int_9_86 bl_int_6_86 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c87
+ bl_int_9_87 bl_int_6_87 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c88
+ bl_int_8_88 wl_0_9 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c0
+ bl_int_10_0 bl_int_8_0 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c1
+ bl_int_10_1 bl_int_8_1 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c2
+ bl_int_8_2 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c3
+ bl_int_8_3 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c4
+ bl_int_10_4 bl_int_9_4 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c5
+ bl_int_10_5 bl_int_9_5 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c6
+ bl_int_9_6 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c7
+ bl_int_9_7 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c8
+ bl_int_10_8 bl_int_8_8 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c9
+ bl_int_10_9 bl_int_8_9 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c10
+ bl_int_8_10 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c11
+ bl_int_8_11 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c12
+ bl_int_10_12 bl_int_9_12 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c13
+ bl_int_10_13 bl_int_9_13 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c14
+ bl_int_9_14 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c15
+ bl_int_9_15 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c16
+ bl_int_10_16 bl_int_8_16 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c17
+ bl_int_10_17 bl_int_8_17 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c18
+ bl_int_8_18 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c19
+ bl_int_8_19 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c20
+ bl_int_10_20 bl_int_9_20 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c21
+ bl_int_10_21 bl_int_9_21 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c22
+ bl_int_9_22 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c23
+ bl_int_9_23 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c24
+ bl_int_10_24 bl_int_8_24 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c25
+ bl_int_10_25 bl_int_8_25 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c26
+ bl_int_8_26 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c27
+ bl_int_8_27 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c28
+ bl_int_10_28 bl_int_9_28 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c29
+ bl_int_10_29 bl_int_9_29 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c30
+ bl_int_9_30 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c31
+ bl_int_9_31 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c32
+ bl_int_10_32 bl_int_8_32 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c33
+ bl_int_10_33 bl_int_8_33 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c34
+ bl_int_8_34 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c35
+ bl_int_8_35 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c36
+ bl_int_10_36 bl_int_9_36 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c37
+ bl_int_10_37 bl_int_9_37 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c38
+ bl_int_9_38 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c39
+ bl_int_9_39 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c40
+ bl_int_10_40 bl_int_8_40 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c41
+ bl_int_10_41 bl_int_8_41 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c42
+ bl_int_8_42 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c43
+ bl_int_8_43 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c44
+ bl_int_10_44 bl_int_9_44 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c45
+ bl_int_10_45 bl_int_9_45 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c46
+ bl_int_9_46 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c47
+ bl_int_9_47 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c48
+ bl_int_10_48 bl_int_8_48 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c49
+ bl_int_10_49 bl_int_8_49 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c50
+ bl_int_8_50 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c51
+ bl_int_8_51 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c52
+ bl_int_10_52 bl_int_9_52 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c53
+ bl_int_10_53 bl_int_9_53 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c54
+ bl_int_9_54 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c55
+ bl_int_9_55 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c56
+ bl_int_10_56 bl_int_8_56 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c57
+ bl_int_10_57 bl_int_8_57 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c58
+ bl_int_8_58 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c59
+ bl_int_8_59 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c60
+ bl_int_10_60 bl_int_9_60 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c61
+ bl_int_10_61 bl_int_9_61 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c62
+ bl_int_9_62 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c63
+ bl_int_9_63 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c64
+ bl_int_10_64 bl_int_8_64 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c65
+ bl_int_10_65 bl_int_8_65 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c66
+ bl_int_8_66 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c67
+ bl_int_8_67 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c68
+ bl_int_10_68 bl_int_9_68 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c69
+ bl_int_10_69 bl_int_9_69 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c70
+ bl_int_9_70 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c71
+ bl_int_9_71 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c72
+ bl_int_10_72 bl_int_8_72 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c73
+ bl_int_10_73 bl_int_8_73 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c74
+ bl_int_8_74 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c75
+ bl_int_8_75 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c76
+ bl_int_10_76 bl_int_9_76 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c77
+ bl_int_10_77 bl_int_9_77 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c78
+ bl_int_9_78 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c79
+ bl_int_9_79 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c80
+ bl_int_10_80 bl_int_8_80 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c81
+ bl_int_10_81 bl_int_8_81 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c82
+ bl_int_8_82 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c83
+ bl_int_8_83 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c84
+ bl_int_10_84 bl_int_9_84 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c85
+ bl_int_10_85 bl_int_9_85 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c86
+ bl_int_9_86 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c87
+ bl_int_9_87 wl_0_10 gnd
+ sram_rom_base_zero_cell
Xbit_r10_c88
+ bl_int_10_88 bl_int_8_88 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r11_c0
+ bl_int_10_0 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c1
+ bl_int_10_1 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c2
+ bl_int_11_2 bl_int_8_2 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c3
+ bl_int_11_3 bl_int_8_3 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c4
+ bl_int_10_4 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c5
+ bl_int_10_5 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c6
+ bl_int_11_6 bl_int_9_6 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c7
+ bl_int_11_7 bl_int_9_7 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c8
+ bl_int_10_8 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c9
+ bl_int_10_9 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c10
+ bl_int_11_10 bl_int_8_10 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c11
+ bl_int_11_11 bl_int_8_11 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c12
+ bl_int_10_12 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c13
+ bl_int_10_13 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c14
+ bl_int_11_14 bl_int_9_14 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c15
+ bl_int_11_15 bl_int_9_15 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c16
+ bl_int_10_16 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c17
+ bl_int_10_17 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c18
+ bl_int_11_18 bl_int_8_18 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c19
+ bl_int_11_19 bl_int_8_19 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c20
+ bl_int_10_20 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c21
+ bl_int_10_21 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c22
+ bl_int_11_22 bl_int_9_22 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c23
+ bl_int_11_23 bl_int_9_23 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c24
+ bl_int_10_24 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c25
+ bl_int_10_25 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c26
+ bl_int_11_26 bl_int_8_26 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c27
+ bl_int_11_27 bl_int_8_27 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c28
+ bl_int_10_28 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c29
+ bl_int_10_29 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c30
+ bl_int_11_30 bl_int_9_30 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c31
+ bl_int_11_31 bl_int_9_31 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c32
+ bl_int_10_32 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c33
+ bl_int_10_33 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c34
+ bl_int_11_34 bl_int_8_34 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c35
+ bl_int_11_35 bl_int_8_35 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c36
+ bl_int_10_36 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c37
+ bl_int_10_37 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c38
+ bl_int_11_38 bl_int_9_38 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c39
+ bl_int_11_39 bl_int_9_39 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c40
+ bl_int_10_40 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c41
+ bl_int_10_41 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c42
+ bl_int_11_42 bl_int_8_42 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c43
+ bl_int_11_43 bl_int_8_43 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c44
+ bl_int_10_44 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c45
+ bl_int_10_45 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c46
+ bl_int_11_46 bl_int_9_46 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c47
+ bl_int_11_47 bl_int_9_47 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c48
+ bl_int_10_48 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c49
+ bl_int_10_49 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c50
+ bl_int_11_50 bl_int_8_50 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c51
+ bl_int_11_51 bl_int_8_51 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c52
+ bl_int_10_52 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c53
+ bl_int_10_53 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c54
+ bl_int_11_54 bl_int_9_54 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c55
+ bl_int_11_55 bl_int_9_55 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c56
+ bl_int_10_56 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c57
+ bl_int_10_57 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c58
+ bl_int_11_58 bl_int_8_58 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c59
+ bl_int_11_59 bl_int_8_59 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c60
+ bl_int_10_60 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c61
+ bl_int_10_61 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c62
+ bl_int_11_62 bl_int_9_62 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c63
+ bl_int_11_63 bl_int_9_63 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c64
+ bl_int_10_64 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c65
+ bl_int_10_65 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c66
+ bl_int_11_66 bl_int_8_66 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c67
+ bl_int_11_67 bl_int_8_67 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c68
+ bl_int_10_68 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c69
+ bl_int_10_69 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c70
+ bl_int_11_70 bl_int_9_70 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c71
+ bl_int_11_71 bl_int_9_71 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c72
+ bl_int_10_72 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c73
+ bl_int_10_73 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c74
+ bl_int_11_74 bl_int_8_74 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c75
+ bl_int_11_75 bl_int_8_75 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c76
+ bl_int_10_76 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c77
+ bl_int_10_77 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c78
+ bl_int_11_78 bl_int_9_78 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c79
+ bl_int_11_79 bl_int_9_79 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c80
+ bl_int_10_80 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c81
+ bl_int_10_81 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c82
+ bl_int_11_82 bl_int_8_82 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c83
+ bl_int_11_83 bl_int_8_83 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c84
+ bl_int_10_84 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c85
+ bl_int_10_85 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r11_c86
+ bl_int_11_86 bl_int_9_86 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c87
+ bl_int_11_87 bl_int_9_87 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c88
+ bl_int_10_88 wl_0_11 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c0
+ bl_int_12_0 bl_int_10_0 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c1
+ bl_int_10_1 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c2
+ bl_int_12_2 bl_int_11_2 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c3
+ bl_int_11_3 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c4
+ bl_int_12_4 bl_int_10_4 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c5
+ bl_int_10_5 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c6
+ bl_int_12_6 bl_int_11_6 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c7
+ bl_int_11_7 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c8
+ bl_int_12_8 bl_int_10_8 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c9
+ bl_int_10_9 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c10
+ bl_int_12_10 bl_int_11_10 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c11
+ bl_int_11_11 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c12
+ bl_int_12_12 bl_int_10_12 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c13
+ bl_int_10_13 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c14
+ bl_int_12_14 bl_int_11_14 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c15
+ bl_int_11_15 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c16
+ bl_int_12_16 bl_int_10_16 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c17
+ bl_int_10_17 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c18
+ bl_int_12_18 bl_int_11_18 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c19
+ bl_int_11_19 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c20
+ bl_int_12_20 bl_int_10_20 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c21
+ bl_int_10_21 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c22
+ bl_int_12_22 bl_int_11_22 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c23
+ bl_int_11_23 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c24
+ bl_int_12_24 bl_int_10_24 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c25
+ bl_int_10_25 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c26
+ bl_int_12_26 bl_int_11_26 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c27
+ bl_int_11_27 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c28
+ bl_int_12_28 bl_int_10_28 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c29
+ bl_int_10_29 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c30
+ bl_int_12_30 bl_int_11_30 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c31
+ bl_int_11_31 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c32
+ bl_int_12_32 bl_int_10_32 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c33
+ bl_int_10_33 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c34
+ bl_int_12_34 bl_int_11_34 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c35
+ bl_int_11_35 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c36
+ bl_int_12_36 bl_int_10_36 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c37
+ bl_int_10_37 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c38
+ bl_int_12_38 bl_int_11_38 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c39
+ bl_int_11_39 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c40
+ bl_int_12_40 bl_int_10_40 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c41
+ bl_int_10_41 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c42
+ bl_int_12_42 bl_int_11_42 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c43
+ bl_int_11_43 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c44
+ bl_int_12_44 bl_int_10_44 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c45
+ bl_int_10_45 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c46
+ bl_int_12_46 bl_int_11_46 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c47
+ bl_int_11_47 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c48
+ bl_int_12_48 bl_int_10_48 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c49
+ bl_int_10_49 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c50
+ bl_int_12_50 bl_int_11_50 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c51
+ bl_int_11_51 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c52
+ bl_int_12_52 bl_int_10_52 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c53
+ bl_int_10_53 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c54
+ bl_int_12_54 bl_int_11_54 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c55
+ bl_int_11_55 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c56
+ bl_int_12_56 bl_int_10_56 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c57
+ bl_int_10_57 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c58
+ bl_int_12_58 bl_int_11_58 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c59
+ bl_int_11_59 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c60
+ bl_int_12_60 bl_int_10_60 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c61
+ bl_int_10_61 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c62
+ bl_int_12_62 bl_int_11_62 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c63
+ bl_int_11_63 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c64
+ bl_int_12_64 bl_int_10_64 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c65
+ bl_int_10_65 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c66
+ bl_int_12_66 bl_int_11_66 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c67
+ bl_int_11_67 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c68
+ bl_int_12_68 bl_int_10_68 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c69
+ bl_int_10_69 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c70
+ bl_int_12_70 bl_int_11_70 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c71
+ bl_int_11_71 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c72
+ bl_int_12_72 bl_int_10_72 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c73
+ bl_int_10_73 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c74
+ bl_int_12_74 bl_int_11_74 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c75
+ bl_int_11_75 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c76
+ bl_int_12_76 bl_int_10_76 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c77
+ bl_int_10_77 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c78
+ bl_int_12_78 bl_int_11_78 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c79
+ bl_int_11_79 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c80
+ bl_int_12_80 bl_int_10_80 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c81
+ bl_int_10_81 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c82
+ bl_int_12_82 bl_int_11_82 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c83
+ bl_int_11_83 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c84
+ bl_int_12_84 bl_int_10_84 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c85
+ bl_int_10_85 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c86
+ bl_int_12_86 bl_int_11_86 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c87
+ bl_int_11_87 wl_0_12 gnd
+ sram_rom_base_zero_cell
Xbit_r12_c88
+ bl_int_12_88 bl_int_10_88 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r13_c0
+ bl_int_12_0 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c1
+ bl_int_13_1 bl_int_10_1 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c2
+ bl_int_12_2 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c3
+ bl_int_13_3 bl_int_11_3 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c4
+ bl_int_12_4 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c5
+ bl_int_13_5 bl_int_10_5 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c6
+ bl_int_12_6 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c7
+ bl_int_13_7 bl_int_11_7 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c8
+ bl_int_12_8 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c9
+ bl_int_13_9 bl_int_10_9 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c10
+ bl_int_12_10 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c11
+ bl_int_13_11 bl_int_11_11 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c12
+ bl_int_12_12 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c13
+ bl_int_13_13 bl_int_10_13 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c14
+ bl_int_12_14 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c15
+ bl_int_13_15 bl_int_11_15 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c16
+ bl_int_12_16 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c17
+ bl_int_13_17 bl_int_10_17 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c18
+ bl_int_12_18 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c19
+ bl_int_13_19 bl_int_11_19 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c20
+ bl_int_12_20 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c21
+ bl_int_13_21 bl_int_10_21 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c22
+ bl_int_12_22 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c23
+ bl_int_13_23 bl_int_11_23 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c24
+ bl_int_12_24 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c25
+ bl_int_13_25 bl_int_10_25 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c26
+ bl_int_12_26 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c27
+ bl_int_13_27 bl_int_11_27 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c28
+ bl_int_12_28 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c29
+ bl_int_13_29 bl_int_10_29 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c30
+ bl_int_12_30 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c31
+ bl_int_13_31 bl_int_11_31 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c32
+ bl_int_12_32 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c33
+ bl_int_13_33 bl_int_10_33 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c34
+ bl_int_12_34 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c35
+ bl_int_13_35 bl_int_11_35 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c36
+ bl_int_12_36 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c37
+ bl_int_13_37 bl_int_10_37 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c38
+ bl_int_12_38 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c39
+ bl_int_13_39 bl_int_11_39 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c40
+ bl_int_12_40 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c41
+ bl_int_13_41 bl_int_10_41 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c42
+ bl_int_12_42 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c43
+ bl_int_13_43 bl_int_11_43 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c44
+ bl_int_12_44 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c45
+ bl_int_13_45 bl_int_10_45 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c46
+ bl_int_12_46 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c47
+ bl_int_13_47 bl_int_11_47 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c48
+ bl_int_12_48 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c49
+ bl_int_13_49 bl_int_10_49 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c50
+ bl_int_12_50 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c51
+ bl_int_13_51 bl_int_11_51 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c52
+ bl_int_12_52 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c53
+ bl_int_13_53 bl_int_10_53 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c54
+ bl_int_12_54 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c55
+ bl_int_13_55 bl_int_11_55 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c56
+ bl_int_12_56 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c57
+ bl_int_13_57 bl_int_10_57 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c58
+ bl_int_12_58 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c59
+ bl_int_13_59 bl_int_11_59 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c60
+ bl_int_12_60 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c61
+ bl_int_13_61 bl_int_10_61 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c62
+ bl_int_12_62 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c63
+ bl_int_13_63 bl_int_11_63 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c64
+ bl_int_12_64 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c65
+ bl_int_13_65 bl_int_10_65 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c66
+ bl_int_12_66 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c67
+ bl_int_13_67 bl_int_11_67 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c68
+ bl_int_12_68 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c69
+ bl_int_13_69 bl_int_10_69 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c70
+ bl_int_12_70 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c71
+ bl_int_13_71 bl_int_11_71 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c72
+ bl_int_12_72 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c73
+ bl_int_13_73 bl_int_10_73 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c74
+ bl_int_12_74 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c75
+ bl_int_13_75 bl_int_11_75 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c76
+ bl_int_12_76 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c77
+ bl_int_13_77 bl_int_10_77 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c78
+ bl_int_12_78 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c79
+ bl_int_13_79 bl_int_11_79 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c80
+ bl_int_12_80 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c81
+ bl_int_13_81 bl_int_10_81 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c82
+ bl_int_12_82 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c83
+ bl_int_13_83 bl_int_11_83 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c84
+ bl_int_12_84 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c85
+ bl_int_13_85 bl_int_10_85 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c86
+ bl_int_12_86 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r13_c87
+ bl_int_13_87 bl_int_11_87 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c88
+ bl_int_12_88 wl_0_13 gnd
+ sram_rom_base_zero_cell
Xbit_r14_c0
+ gnd bl_int_12_0 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c1
+ gnd bl_int_13_1 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c2
+ gnd bl_int_12_2 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c3
+ gnd bl_int_13_3 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c4
+ gnd bl_int_12_4 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c5
+ gnd bl_int_13_5 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c6
+ gnd bl_int_12_6 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c7
+ gnd bl_int_13_7 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c8
+ gnd bl_int_12_8 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c9
+ gnd bl_int_13_9 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c10
+ gnd bl_int_12_10 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c11
+ gnd bl_int_13_11 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c12
+ gnd bl_int_12_12 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c13
+ gnd bl_int_13_13 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c14
+ gnd bl_int_12_14 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c15
+ gnd bl_int_13_15 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c16
+ gnd bl_int_12_16 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c17
+ gnd bl_int_13_17 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c18
+ gnd bl_int_12_18 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c19
+ gnd bl_int_13_19 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c20
+ gnd bl_int_12_20 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c21
+ gnd bl_int_13_21 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c22
+ gnd bl_int_12_22 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c23
+ gnd bl_int_13_23 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c24
+ gnd bl_int_12_24 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c25
+ gnd bl_int_13_25 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c26
+ gnd bl_int_12_26 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c27
+ gnd bl_int_13_27 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c28
+ gnd bl_int_12_28 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c29
+ gnd bl_int_13_29 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c30
+ gnd bl_int_12_30 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c31
+ gnd bl_int_13_31 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c32
+ gnd bl_int_12_32 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c33
+ gnd bl_int_13_33 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c34
+ gnd bl_int_12_34 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c35
+ gnd bl_int_13_35 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c36
+ gnd bl_int_12_36 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c37
+ gnd bl_int_13_37 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c38
+ gnd bl_int_12_38 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c39
+ gnd bl_int_13_39 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c40
+ gnd bl_int_12_40 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c41
+ gnd bl_int_13_41 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c42
+ gnd bl_int_12_42 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c43
+ gnd bl_int_13_43 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c44
+ gnd bl_int_12_44 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c45
+ gnd bl_int_13_45 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c46
+ gnd bl_int_12_46 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c47
+ gnd bl_int_13_47 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c48
+ gnd bl_int_12_48 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c49
+ gnd bl_int_13_49 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c50
+ gnd bl_int_12_50 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c51
+ gnd bl_int_13_51 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c52
+ gnd bl_int_12_52 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c53
+ gnd bl_int_13_53 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c54
+ gnd bl_int_12_54 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c55
+ gnd bl_int_13_55 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c56
+ gnd bl_int_12_56 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c57
+ gnd bl_int_13_57 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c58
+ gnd bl_int_12_58 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c59
+ gnd bl_int_13_59 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c60
+ gnd bl_int_12_60 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c61
+ gnd bl_int_13_61 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c62
+ gnd bl_int_12_62 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c63
+ gnd bl_int_13_63 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c64
+ gnd bl_int_12_64 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c65
+ gnd bl_int_13_65 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c66
+ gnd bl_int_12_66 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c67
+ gnd bl_int_13_67 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c68
+ gnd bl_int_12_68 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c69
+ gnd bl_int_13_69 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c70
+ gnd bl_int_12_70 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c71
+ gnd bl_int_13_71 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c72
+ gnd bl_int_12_72 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c73
+ gnd bl_int_13_73 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c74
+ gnd bl_int_12_74 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c75
+ gnd bl_int_13_75 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c76
+ gnd bl_int_12_76 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c77
+ gnd bl_int_13_77 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c78
+ gnd bl_int_12_78 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c79
+ gnd bl_int_13_79 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c80
+ gnd bl_int_12_80 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c81
+ gnd bl_int_13_81 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c82
+ gnd bl_int_12_82 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c83
+ gnd bl_int_13_83 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c84
+ gnd bl_int_12_84 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c85
+ gnd bl_int_13_85 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c86
+ gnd bl_int_12_86 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c87
+ gnd bl_int_13_87 precharge gnd
+ sram_rom_base_one_cell
Xbit_r14_c88
+ gnd bl_int_12_88 precharge gnd
+ sram_rom_base_one_cell
Xbitcell_array_precharge
+ bl_0_0 bl_0_1 bl_0_2 bl_0_3 bl_0_4 bl_0_5 bl_0_6 bl_0_7 bl_0_8 bl_0_9
+ bl_0_10 bl_0_11 bl_0_12 bl_0_13 bl_0_14 bl_0_15 bl_0_16 bl_0_17
+ bl_0_18 bl_0_19 bl_0_20 bl_0_21 bl_0_22 bl_0_23 bl_0_24 bl_0_25
+ bl_0_26 bl_0_27 bl_0_28 bl_0_29 bl_0_30 bl_0_31 bl_0_32 bl_0_33
+ bl_0_34 bl_0_35 bl_0_36 bl_0_37 bl_0_38 bl_0_39 bl_0_40 bl_0_41
+ bl_0_42 bl_0_43 bl_0_44 bl_0_45 bl_0_46 bl_0_47 bl_0_48 bl_0_49
+ bl_0_50 bl_0_51 bl_0_52 bl_0_53 bl_0_54 bl_0_55 bl_0_56 bl_0_57
+ bl_0_58 bl_0_59 bl_0_60 bl_0_61 bl_0_62 bl_0_63 bl_0_64 bl_0_65
+ bl_0_66 bl_0_67 bl_0_68 bl_0_69 bl_0_70 bl_0_71 bl_0_72 bl_0_73
+ bl_0_74 bl_0_75 bl_0_76 bl_0_77 bl_0_78 bl_0_79 bl_0_80 bl_0_81
+ bl_0_82 bl_0_83 bl_0_84 bl_0_85 bl_0_86 bl_0_87 bl_0_88 precharge vdd
+ sram_rom_precharge_array_0
.ENDS sram_rom_row_decode_array

.SUBCKT sram_rom_address_control_array
+ A0_in A1_in A2_in A3_in A4_in A5_in A6_in A0_out A1_out A2_out A3_out
+ A4_out A5_out A6_out Abar0_out Abar1_out Abar2_out Abar3_out Abar4_out
+ Abar5_out Abar6_out clk vdd gnd
* INPUT : A0_in 
* INPUT : A1_in 
* INPUT : A2_in 
* INPUT : A3_in 
* INPUT : A4_in 
* INPUT : A5_in 
* INPUT : A6_in 
* OUTPUT: A0_out 
* OUTPUT: A1_out 
* OUTPUT: A2_out 
* OUTPUT: A3_out 
* OUTPUT: A4_out 
* OUTPUT: A5_out 
* OUTPUT: A6_out 
* OUTPUT: Abar0_out 
* OUTPUT: Abar1_out 
* OUTPUT: Abar2_out 
* OUTPUT: Abar3_out 
* OUTPUT: Abar4_out 
* OUTPUT: Abar5_out 
* OUTPUT: Abar6_out 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
XXaddr_buf_0
+ A0_in A0_out Abar0_out clk vdd gnd
+ sram_rom_address_control_buf
XXaddr_buf_1
+ A1_in A1_out Abar1_out clk vdd gnd
+ sram_rom_address_control_buf
XXaddr_buf_2
+ A2_in A2_out Abar2_out clk vdd gnd
+ sram_rom_address_control_buf
XXaddr_buf_3
+ A3_in A3_out Abar3_out clk vdd gnd
+ sram_rom_address_control_buf
XXaddr_buf_4
+ A4_in A4_out Abar4_out clk vdd gnd
+ sram_rom_address_control_buf
XXaddr_buf_5
+ A5_in A5_out Abar5_out clk vdd gnd
+ sram_rom_address_control_buf
XXaddr_buf_6
+ A6_in A6_out Abar6_out clk vdd gnd
+ sram_rom_address_control_buf
.ENDS sram_rom_address_control_array

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u

.SUBCKT sram_pinv_dec_1
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
.ENDS sram_pinv_dec_1

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT sram_pinv_dec_0
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS sram_pinv_dec_0

.SUBCKT sram_pbuf_dec
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xbuf_inv1
+ A zb_int vdd gnd
+ sram_pinv_dec_0
Xbuf_inv2
+ zb_int Z vdd gnd
+ sram_pinv_dec_1
.ENDS sram_pbuf_dec

.SUBCKT sram_rom_row_decode_wordline_buffer
+ in_0 in_1 in_2 in_3 in_4 in_5 in_6 in_7 in_8 in_9 in_10 in_11 in_12
+ in_13 in_14 in_15 in_16 in_17 in_18 in_19 in_20 in_21 in_22 in_23
+ in_24 in_25 in_26 in_27 in_28 in_29 in_30 in_31 in_32 in_33 in_34
+ in_35 in_36 in_37 in_38 in_39 in_40 in_41 in_42 in_43 in_44 in_45
+ in_46 in_47 in_48 in_49 in_50 in_51 in_52 in_53 in_54 in_55 in_56
+ in_57 in_58 in_59 in_60 in_61 in_62 in_63 in_64 in_65 in_66 in_67
+ in_68 in_69 in_70 in_71 in_72 in_73 in_74 in_75 in_76 in_77 in_78
+ in_79 in_80 in_81 in_82 in_83 in_84 in_85 in_86 in_87 in_88 out_0
+ out_1 out_2 out_3 out_4 out_5 out_6 out_7 out_8 out_9 out_10 out_11
+ out_12 out_13 out_14 out_15 out_16 out_17 out_18 out_19 out_20 out_21
+ out_22 out_23 out_24 out_25 out_26 out_27 out_28 out_29 out_30 out_31
+ out_32 out_33 out_34 out_35 out_36 out_37 out_38 out_39 out_40 out_41
+ out_42 out_43 out_44 out_45 out_46 out_47 out_48 out_49 out_50 out_51
+ out_52 out_53 out_54 out_55 out_56 out_57 out_58 out_59 out_60 out_61
+ out_62 out_63 out_64 out_65 out_66 out_67 out_68 out_69 out_70 out_71
+ out_72 out_73 out_74 out_75 out_76 out_77 out_78 out_79 out_80 out_81
+ out_82 out_83 out_84 out_85 out_86 out_87 out_88 vdd gnd
* INPUT : in_0 
* INPUT : in_1 
* INPUT : in_2 
* INPUT : in_3 
* INPUT : in_4 
* INPUT : in_5 
* INPUT : in_6 
* INPUT : in_7 
* INPUT : in_8 
* INPUT : in_9 
* INPUT : in_10 
* INPUT : in_11 
* INPUT : in_12 
* INPUT : in_13 
* INPUT : in_14 
* INPUT : in_15 
* INPUT : in_16 
* INPUT : in_17 
* INPUT : in_18 
* INPUT : in_19 
* INPUT : in_20 
* INPUT : in_21 
* INPUT : in_22 
* INPUT : in_23 
* INPUT : in_24 
* INPUT : in_25 
* INPUT : in_26 
* INPUT : in_27 
* INPUT : in_28 
* INPUT : in_29 
* INPUT : in_30 
* INPUT : in_31 
* INPUT : in_32 
* INPUT : in_33 
* INPUT : in_34 
* INPUT : in_35 
* INPUT : in_36 
* INPUT : in_37 
* INPUT : in_38 
* INPUT : in_39 
* INPUT : in_40 
* INPUT : in_41 
* INPUT : in_42 
* INPUT : in_43 
* INPUT : in_44 
* INPUT : in_45 
* INPUT : in_46 
* INPUT : in_47 
* INPUT : in_48 
* INPUT : in_49 
* INPUT : in_50 
* INPUT : in_51 
* INPUT : in_52 
* INPUT : in_53 
* INPUT : in_54 
* INPUT : in_55 
* INPUT : in_56 
* INPUT : in_57 
* INPUT : in_58 
* INPUT : in_59 
* INPUT : in_60 
* INPUT : in_61 
* INPUT : in_62 
* INPUT : in_63 
* INPUT : in_64 
* INPUT : in_65 
* INPUT : in_66 
* INPUT : in_67 
* INPUT : in_68 
* INPUT : in_69 
* INPUT : in_70 
* INPUT : in_71 
* INPUT : in_72 
* INPUT : in_73 
* INPUT : in_74 
* INPUT : in_75 
* INPUT : in_76 
* INPUT : in_77 
* INPUT : in_78 
* INPUT : in_79 
* INPUT : in_80 
* INPUT : in_81 
* INPUT : in_82 
* INPUT : in_83 
* INPUT : in_84 
* INPUT : in_85 
* INPUT : in_86 
* INPUT : in_87 
* INPUT : in_88 
* OUTPUT: out_0 
* OUTPUT: out_1 
* OUTPUT: out_2 
* OUTPUT: out_3 
* OUTPUT: out_4 
* OUTPUT: out_5 
* OUTPUT: out_6 
* OUTPUT: out_7 
* OUTPUT: out_8 
* OUTPUT: out_9 
* OUTPUT: out_10 
* OUTPUT: out_11 
* OUTPUT: out_12 
* OUTPUT: out_13 
* OUTPUT: out_14 
* OUTPUT: out_15 
* OUTPUT: out_16 
* OUTPUT: out_17 
* OUTPUT: out_18 
* OUTPUT: out_19 
* OUTPUT: out_20 
* OUTPUT: out_21 
* OUTPUT: out_22 
* OUTPUT: out_23 
* OUTPUT: out_24 
* OUTPUT: out_25 
* OUTPUT: out_26 
* OUTPUT: out_27 
* OUTPUT: out_28 
* OUTPUT: out_29 
* OUTPUT: out_30 
* OUTPUT: out_31 
* OUTPUT: out_32 
* OUTPUT: out_33 
* OUTPUT: out_34 
* OUTPUT: out_35 
* OUTPUT: out_36 
* OUTPUT: out_37 
* OUTPUT: out_38 
* OUTPUT: out_39 
* OUTPUT: out_40 
* OUTPUT: out_41 
* OUTPUT: out_42 
* OUTPUT: out_43 
* OUTPUT: out_44 
* OUTPUT: out_45 
* OUTPUT: out_46 
* OUTPUT: out_47 
* OUTPUT: out_48 
* OUTPUT: out_49 
* OUTPUT: out_50 
* OUTPUT: out_51 
* OUTPUT: out_52 
* OUTPUT: out_53 
* OUTPUT: out_54 
* OUTPUT: out_55 
* OUTPUT: out_56 
* OUTPUT: out_57 
* OUTPUT: out_58 
* OUTPUT: out_59 
* OUTPUT: out_60 
* OUTPUT: out_61 
* OUTPUT: out_62 
* OUTPUT: out_63 
* OUTPUT: out_64 
* OUTPUT: out_65 
* OUTPUT: out_66 
* OUTPUT: out_67 
* OUTPUT: out_68 
* OUTPUT: out_69 
* OUTPUT: out_70 
* OUTPUT: out_71 
* OUTPUT: out_72 
* OUTPUT: out_73 
* OUTPUT: out_74 
* OUTPUT: out_75 
* OUTPUT: out_76 
* OUTPUT: out_77 
* OUTPUT: out_78 
* OUTPUT: out_79 
* OUTPUT: out_80 
* OUTPUT: out_81 
* OUTPUT: out_82 
* OUTPUT: out_83 
* OUTPUT: out_84 
* OUTPUT: out_85 
* OUTPUT: out_86 
* OUTPUT: out_87 
* OUTPUT: out_88 
* POWER : vdd 
* GROUND: gnd 
* rows: 89 Buffer size of: 23
Xwld0
+ in_0 out_0 vdd gnd
+ sram_pbuf_dec
Xwld1
+ in_1 out_1 vdd gnd
+ sram_pbuf_dec
Xwld2
+ in_2 out_2 vdd gnd
+ sram_pbuf_dec
Xwld3
+ in_3 out_3 vdd gnd
+ sram_pbuf_dec
Xwld4
+ in_4 out_4 vdd gnd
+ sram_pbuf_dec
Xwld5
+ in_5 out_5 vdd gnd
+ sram_pbuf_dec
Xwld6
+ in_6 out_6 vdd gnd
+ sram_pbuf_dec
Xwld7
+ in_7 out_7 vdd gnd
+ sram_pbuf_dec
Xwld8
+ in_8 out_8 vdd gnd
+ sram_pbuf_dec
Xwld9
+ in_9 out_9 vdd gnd
+ sram_pbuf_dec
Xwld10
+ in_10 out_10 vdd gnd
+ sram_pbuf_dec
Xwld11
+ in_11 out_11 vdd gnd
+ sram_pbuf_dec
Xwld12
+ in_12 out_12 vdd gnd
+ sram_pbuf_dec
Xwld13
+ in_13 out_13 vdd gnd
+ sram_pbuf_dec
Xwld14
+ in_14 out_14 vdd gnd
+ sram_pbuf_dec
Xwld15
+ in_15 out_15 vdd gnd
+ sram_pbuf_dec
Xwld16
+ in_16 out_16 vdd gnd
+ sram_pbuf_dec
Xwld17
+ in_17 out_17 vdd gnd
+ sram_pbuf_dec
Xwld18
+ in_18 out_18 vdd gnd
+ sram_pbuf_dec
Xwld19
+ in_19 out_19 vdd gnd
+ sram_pbuf_dec
Xwld20
+ in_20 out_20 vdd gnd
+ sram_pbuf_dec
Xwld21
+ in_21 out_21 vdd gnd
+ sram_pbuf_dec
Xwld22
+ in_22 out_22 vdd gnd
+ sram_pbuf_dec
Xwld23
+ in_23 out_23 vdd gnd
+ sram_pbuf_dec
Xwld24
+ in_24 out_24 vdd gnd
+ sram_pbuf_dec
Xwld25
+ in_25 out_25 vdd gnd
+ sram_pbuf_dec
Xwld26
+ in_26 out_26 vdd gnd
+ sram_pbuf_dec
Xwld27
+ in_27 out_27 vdd gnd
+ sram_pbuf_dec
Xwld28
+ in_28 out_28 vdd gnd
+ sram_pbuf_dec
Xwld29
+ in_29 out_29 vdd gnd
+ sram_pbuf_dec
Xwld30
+ in_30 out_30 vdd gnd
+ sram_pbuf_dec
Xwld31
+ in_31 out_31 vdd gnd
+ sram_pbuf_dec
Xwld32
+ in_32 out_32 vdd gnd
+ sram_pbuf_dec
Xwld33
+ in_33 out_33 vdd gnd
+ sram_pbuf_dec
Xwld34
+ in_34 out_34 vdd gnd
+ sram_pbuf_dec
Xwld35
+ in_35 out_35 vdd gnd
+ sram_pbuf_dec
Xwld36
+ in_36 out_36 vdd gnd
+ sram_pbuf_dec
Xwld37
+ in_37 out_37 vdd gnd
+ sram_pbuf_dec
Xwld38
+ in_38 out_38 vdd gnd
+ sram_pbuf_dec
Xwld39
+ in_39 out_39 vdd gnd
+ sram_pbuf_dec
Xwld40
+ in_40 out_40 vdd gnd
+ sram_pbuf_dec
Xwld41
+ in_41 out_41 vdd gnd
+ sram_pbuf_dec
Xwld42
+ in_42 out_42 vdd gnd
+ sram_pbuf_dec
Xwld43
+ in_43 out_43 vdd gnd
+ sram_pbuf_dec
Xwld44
+ in_44 out_44 vdd gnd
+ sram_pbuf_dec
Xwld45
+ in_45 out_45 vdd gnd
+ sram_pbuf_dec
Xwld46
+ in_46 out_46 vdd gnd
+ sram_pbuf_dec
Xwld47
+ in_47 out_47 vdd gnd
+ sram_pbuf_dec
Xwld48
+ in_48 out_48 vdd gnd
+ sram_pbuf_dec
Xwld49
+ in_49 out_49 vdd gnd
+ sram_pbuf_dec
Xwld50
+ in_50 out_50 vdd gnd
+ sram_pbuf_dec
Xwld51
+ in_51 out_51 vdd gnd
+ sram_pbuf_dec
Xwld52
+ in_52 out_52 vdd gnd
+ sram_pbuf_dec
Xwld53
+ in_53 out_53 vdd gnd
+ sram_pbuf_dec
Xwld54
+ in_54 out_54 vdd gnd
+ sram_pbuf_dec
Xwld55
+ in_55 out_55 vdd gnd
+ sram_pbuf_dec
Xwld56
+ in_56 out_56 vdd gnd
+ sram_pbuf_dec
Xwld57
+ in_57 out_57 vdd gnd
+ sram_pbuf_dec
Xwld58
+ in_58 out_58 vdd gnd
+ sram_pbuf_dec
Xwld59
+ in_59 out_59 vdd gnd
+ sram_pbuf_dec
Xwld60
+ in_60 out_60 vdd gnd
+ sram_pbuf_dec
Xwld61
+ in_61 out_61 vdd gnd
+ sram_pbuf_dec
Xwld62
+ in_62 out_62 vdd gnd
+ sram_pbuf_dec
Xwld63
+ in_63 out_63 vdd gnd
+ sram_pbuf_dec
Xwld64
+ in_64 out_64 vdd gnd
+ sram_pbuf_dec
Xwld65
+ in_65 out_65 vdd gnd
+ sram_pbuf_dec
Xwld66
+ in_66 out_66 vdd gnd
+ sram_pbuf_dec
Xwld67
+ in_67 out_67 vdd gnd
+ sram_pbuf_dec
Xwld68
+ in_68 out_68 vdd gnd
+ sram_pbuf_dec
Xwld69
+ in_69 out_69 vdd gnd
+ sram_pbuf_dec
Xwld70
+ in_70 out_70 vdd gnd
+ sram_pbuf_dec
Xwld71
+ in_71 out_71 vdd gnd
+ sram_pbuf_dec
Xwld72
+ in_72 out_72 vdd gnd
+ sram_pbuf_dec
Xwld73
+ in_73 out_73 vdd gnd
+ sram_pbuf_dec
Xwld74
+ in_74 out_74 vdd gnd
+ sram_pbuf_dec
Xwld75
+ in_75 out_75 vdd gnd
+ sram_pbuf_dec
Xwld76
+ in_76 out_76 vdd gnd
+ sram_pbuf_dec
Xwld77
+ in_77 out_77 vdd gnd
+ sram_pbuf_dec
Xwld78
+ in_78 out_78 vdd gnd
+ sram_pbuf_dec
Xwld79
+ in_79 out_79 vdd gnd
+ sram_pbuf_dec
Xwld80
+ in_80 out_80 vdd gnd
+ sram_pbuf_dec
Xwld81
+ in_81 out_81 vdd gnd
+ sram_pbuf_dec
Xwld82
+ in_82 out_82 vdd gnd
+ sram_pbuf_dec
Xwld83
+ in_83 out_83 vdd gnd
+ sram_pbuf_dec
Xwld84
+ in_84 out_84 vdd gnd
+ sram_pbuf_dec
Xwld85
+ in_85 out_85 vdd gnd
+ sram_pbuf_dec
Xwld86
+ in_86 out_86 vdd gnd
+ sram_pbuf_dec
Xwld87
+ in_87 out_87 vdd gnd
+ sram_pbuf_dec
Xwld88
+ in_88 out_88 vdd gnd
+ sram_pbuf_dec
.ENDS sram_rom_row_decode_wordline_buffer

.SUBCKT sram_rom_row_decode
+ A0 A1 A2 A3 A4 A5 A6 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9
+ wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20
+ wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31
+ wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42
+ wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53
+ wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64
+ wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75
+ wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86
+ wl_87 wl_88 precharge clk vdd gnd
* INPUT : A0 
* INPUT : A1 
* INPUT : A2 
* INPUT : A3 
* INPUT : A4 
* INPUT : A5 
* INPUT : A6 
* OUTPUT: wl_0 
* OUTPUT: wl_1 
* OUTPUT: wl_2 
* OUTPUT: wl_3 
* OUTPUT: wl_4 
* OUTPUT: wl_5 
* OUTPUT: wl_6 
* OUTPUT: wl_7 
* OUTPUT: wl_8 
* OUTPUT: wl_9 
* OUTPUT: wl_10 
* OUTPUT: wl_11 
* OUTPUT: wl_12 
* OUTPUT: wl_13 
* OUTPUT: wl_14 
* OUTPUT: wl_15 
* OUTPUT: wl_16 
* OUTPUT: wl_17 
* OUTPUT: wl_18 
* OUTPUT: wl_19 
* OUTPUT: wl_20 
* OUTPUT: wl_21 
* OUTPUT: wl_22 
* OUTPUT: wl_23 
* OUTPUT: wl_24 
* OUTPUT: wl_25 
* OUTPUT: wl_26 
* OUTPUT: wl_27 
* OUTPUT: wl_28 
* OUTPUT: wl_29 
* OUTPUT: wl_30 
* OUTPUT: wl_31 
* OUTPUT: wl_32 
* OUTPUT: wl_33 
* OUTPUT: wl_34 
* OUTPUT: wl_35 
* OUTPUT: wl_36 
* OUTPUT: wl_37 
* OUTPUT: wl_38 
* OUTPUT: wl_39 
* OUTPUT: wl_40 
* OUTPUT: wl_41 
* OUTPUT: wl_42 
* OUTPUT: wl_43 
* OUTPUT: wl_44 
* OUTPUT: wl_45 
* OUTPUT: wl_46 
* OUTPUT: wl_47 
* OUTPUT: wl_48 
* OUTPUT: wl_49 
* OUTPUT: wl_50 
* OUTPUT: wl_51 
* OUTPUT: wl_52 
* OUTPUT: wl_53 
* OUTPUT: wl_54 
* OUTPUT: wl_55 
* OUTPUT: wl_56 
* OUTPUT: wl_57 
* OUTPUT: wl_58 
* OUTPUT: wl_59 
* OUTPUT: wl_60 
* OUTPUT: wl_61 
* OUTPUT: wl_62 
* OUTPUT: wl_63 
* OUTPUT: wl_64 
* OUTPUT: wl_65 
* OUTPUT: wl_66 
* OUTPUT: wl_67 
* OUTPUT: wl_68 
* OUTPUT: wl_69 
* OUTPUT: wl_70 
* OUTPUT: wl_71 
* OUTPUT: wl_72 
* OUTPUT: wl_73 
* OUTPUT: wl_74 
* OUTPUT: wl_75 
* OUTPUT: wl_76 
* OUTPUT: wl_77 
* OUTPUT: wl_78 
* OUTPUT: wl_79 
* OUTPUT: wl_80 
* OUTPUT: wl_81 
* OUTPUT: wl_82 
* OUTPUT: wl_83 
* OUTPUT: wl_84 
* OUTPUT: wl_85 
* OUTPUT: wl_86 
* OUTPUT: wl_87 
* OUTPUT: wl_88 
* INPUT : precharge 
* INPUT : clk 
* POWER : vdd 
* GROUND: gnd 
Xdecode_array_inst
+ wl_int0 wl_int1 wl_int2 wl_int3 wl_int4 wl_int5 wl_int6 wl_int7
+ wl_int8 wl_int9 wl_int10 wl_int11 wl_int12 wl_int13 wl_int14 wl_int15
+ wl_int16 wl_int17 wl_int18 wl_int19 wl_int20 wl_int21 wl_int22
+ wl_int23 wl_int24 wl_int25 wl_int26 wl_int27 wl_int28 wl_int29
+ wl_int30 wl_int31 wl_int32 wl_int33 wl_int34 wl_int35 wl_int36
+ wl_int37 wl_int38 wl_int39 wl_int40 wl_int41 wl_int42 wl_int43
+ wl_int44 wl_int45 wl_int46 wl_int47 wl_int48 wl_int49 wl_int50
+ wl_int51 wl_int52 wl_int53 wl_int54 wl_int55 wl_int56 wl_int57
+ wl_int58 wl_int59 wl_int60 wl_int61 wl_int62 wl_int63 wl_int64
+ wl_int65 wl_int66 wl_int67 wl_int68 wl_int69 wl_int70 wl_int71
+ wl_int72 wl_int73 wl_int74 wl_int75 wl_int76 wl_int77 wl_int78
+ wl_int79 wl_int80 wl_int81 wl_int82 wl_int83 wl_int84 wl_int85
+ wl_int86 wl_int87 wl_int88 Ab_int_6 A_int_6 Ab_int_5 A_int_5 Ab_int_4
+ A_int_4 Ab_int_3 A_int_3 Ab_int_2 A_int_2 Ab_int_1 A_int_1 Ab_int_0
+ A_int_0 precharge vdd gnd
+ sram_rom_row_decode_array
Xpre_control_array
+ A0 A1 A2 A3 A4 A5 A6 A_int_0 A_int_1 A_int_2 A_int_3 A_int_4 A_int_5
+ A_int_6 Ab_int_0 Ab_int_1 Ab_int_2 Ab_int_3 Ab_int_4 Ab_int_5 Ab_int_6
+ clk vdd gnd
+ sram_rom_address_control_array
Xrom_wordline_driver
+ wl_int0 wl_int1 wl_int2 wl_int3 wl_int4 wl_int5 wl_int6 wl_int7
+ wl_int8 wl_int9 wl_int10 wl_int11 wl_int12 wl_int13 wl_int14 wl_int15
+ wl_int16 wl_int17 wl_int18 wl_int19 wl_int20 wl_int21 wl_int22
+ wl_int23 wl_int24 wl_int25 wl_int26 wl_int27 wl_int28 wl_int29
+ wl_int30 wl_int31 wl_int32 wl_int33 wl_int34 wl_int35 wl_int36
+ wl_int37 wl_int38 wl_int39 wl_int40 wl_int41 wl_int42 wl_int43
+ wl_int44 wl_int45 wl_int46 wl_int47 wl_int48 wl_int49 wl_int50
+ wl_int51 wl_int52 wl_int53 wl_int54 wl_int55 wl_int56 wl_int57
+ wl_int58 wl_int59 wl_int60 wl_int61 wl_int62 wl_int63 wl_int64
+ wl_int65 wl_int66 wl_int67 wl_int68 wl_int69 wl_int70 wl_int71
+ wl_int72 wl_int73 wl_int74 wl_int75 wl_int76 wl_int77 wl_int78
+ wl_int79 wl_int80 wl_int81 wl_int82 wl_int83 wl_int84 wl_int85
+ wl_int86 wl_int87 wl_int88 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7
+ wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19
+ wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30
+ wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41
+ wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52
+ wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63
+ wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74
+ wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85
+ wl_86 wl_87 wl_88 vdd gnd
+ sram_rom_row_decode_wordline_buffer
.ENDS sram_rom_row_decode

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=4 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=4 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT sram_pinv_1
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=4 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=4 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
.ENDS sram_pinv_1

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=2 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u

.SUBCKT sram_pinv_0
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=2 w=2.0 l=0.15 pd=4.30 ps=4.30 as=0.75u ad=0.75u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=2 w=1.26 l=0.15 pd=2.82 ps=2.82 as=0.47u ad=0.47u
.ENDS sram_pinv_0

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u

.SUBCKT sram_pinv
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.36 l=0.15 pd=1.02 ps=1.02 as=0.14u ad=0.14u
.ENDS sram_pinv

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=7 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=7 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

.SUBCKT sram_pinv_2
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=7 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=7 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u
.ENDS sram_pinv_2

.SUBCKT sram_rom_clock_driver
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 1, 3, 10, 31]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ sram_pinv
Xbuf_inv2
+ Zb1_int Zb2_int vdd gnd
+ sram_pinv
Xbuf_inv3
+ Zb2_int Zb3_int vdd gnd
+ sram_pinv
Xbuf_inv4
+ Zb3_int Zb4_int vdd gnd
+ sram_pinv_0
Xbuf_inv5
+ Zb4_int Zb5_int vdd gnd
+ sram_pinv_1
Xbuf_inv6
+ Zb5_int Z vdd gnd
+ sram_pinv_2
.ENDS sram_rom_clock_driver

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=16 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=16 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

.SUBCKT sram_pinv_5
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=16 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=16 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
.ENDS sram_pinv_5

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u

.SUBCKT sram_pinv_3
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=3.0 l=0.15 pd=6.30 ps=6.30 as=1.12u ad=1.12u
.ENDS sram_pinv_3

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=6 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=6 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u

.SUBCKT sram_pinv_4
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpinv_pmos Z A vdd vdd sky130_fd_pr__pfet_01v8 m=6 w=5.0 l=0.15 pd=10.30 ps=10.30 as=1.88u ad=1.88u
Xpinv_nmos Z A gnd gnd sky130_fd_pr__nfet_01v8 m=6 w=7.0 l=0.15 pd=14.30 ps=14.30 as=2.62u ad=2.62u
.ENDS sram_pinv_4

.SUBCKT sram_rom_precharge_driver
+ A Z vdd gnd
* INPUT : A 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
* sizes: [1, 1, 1, 3, 8, 24, 73]
Xbuf_inv1
+ A Zb1_int vdd gnd
+ sram_pinv
Xbuf_inv2
+ Zb1_int Zb2_int vdd gnd
+ sram_pinv
Xbuf_inv3
+ Zb2_int Zb3_int vdd gnd
+ sram_pinv
Xbuf_inv4
+ Zb3_int Zb4_int vdd gnd
+ sram_pinv_0
Xbuf_inv5
+ Zb4_int Zb5_int vdd gnd
+ sram_pinv_3
Xbuf_inv6
+ Zb5_int Zb6_int vdd gnd
+ sram_pinv_4
Xbuf_inv7
+ Zb6_int Z vdd gnd
+ sram_pinv_5
.ENDS sram_rom_precharge_driver

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

* spice ptx X{0} {1} sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u

* spice ptx X{0} {1} sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u

.SUBCKT sram_rom_control_nand
+ A B Z vdd gnd
* INPUT : A 
* INPUT : B 
* OUTPUT: Z 
* POWER : vdd 
* GROUND: gnd 
Xpnand2_pmos1 vdd A Z vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_pmos2 Z B vdd vdd sky130_fd_pr__pfet_01v8 m=1 w=1.12 l=0.15 pd=2.54 ps=2.54 as=0.42u ad=0.42u
Xpnand2_nmos1 Z B net1 gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
Xpnand2_nmos2 net1 A gnd gnd sky130_fd_pr__nfet_01v8 m=1 w=0.74 l=0.15 pd=1.78 ps=1.78 as=0.28u ad=0.28u
.ENDS sram_rom_control_nand

.SUBCKT sram_rom_control_logic
+ clk_in CS prechrg clk_out vdd gnd
* INPUT : clk_in 
* INPUT : CS 
* OUTPUT: prechrg 
* OUTPUT: clk_out 
* POWER : vdd 
* GROUND: gnd 
Xclk_driver
+ clk_in clk_out vdd gnd
+ sram_rom_clock_driver
Xcontrol_nand
+ CS clk_out pre_drive vdd gnd
+ sram_rom_control_nand
Xprecharge_driver
+ pre_drive prechrg vdd gnd
+ sram_rom_precharge_driver
.ENDS sram_rom_control_logic

.SUBCKT sram_rom_precharge_array
+ pre_bl0_out pre_bl1_out pre_bl2_out pre_bl3_out pre_bl4_out
+ pre_bl5_out pre_bl6_out pre_bl7_out pre_bl8_out pre_bl9_out
+ pre_bl10_out pre_bl11_out pre_bl12_out pre_bl13_out pre_bl14_out
+ pre_bl15_out pre_bl16_out pre_bl17_out pre_bl18_out pre_bl19_out
+ pre_bl20_out pre_bl21_out pre_bl22_out pre_bl23_out pre_bl24_out
+ pre_bl25_out pre_bl26_out pre_bl27_out pre_bl28_out pre_bl29_out
+ pre_bl30_out pre_bl31_out pre_bl32_out pre_bl33_out pre_bl34_out
+ pre_bl35_out pre_bl36_out pre_bl37_out pre_bl38_out pre_bl39_out
+ pre_bl40_out pre_bl41_out pre_bl42_out pre_bl43_out pre_bl44_out
+ pre_bl45_out pre_bl46_out pre_bl47_out pre_bl48_out pre_bl49_out
+ pre_bl50_out pre_bl51_out pre_bl52_out pre_bl53_out pre_bl54_out
+ pre_bl55_out pre_bl56_out pre_bl57_out pre_bl58_out pre_bl59_out
+ pre_bl60_out pre_bl61_out pre_bl62_out pre_bl63_out pre_bl64_out
+ pre_bl65_out pre_bl66_out pre_bl67_out pre_bl68_out pre_bl69_out
+ pre_bl70_out pre_bl71_out pre_bl72_out pre_bl73_out pre_bl74_out
+ pre_bl75_out pre_bl76_out pre_bl77_out pre_bl78_out pre_bl79_out
+ pre_bl80_out pre_bl81_out pre_bl82_out pre_bl83_out pre_bl84_out
+ pre_bl85_out pre_bl86_out pre_bl87_out pre_bl88_out pre_bl89_out
+ pre_bl90_out pre_bl91_out pre_bl92_out pre_bl93_out pre_bl94_out
+ pre_bl95_out pre_bl96_out pre_bl97_out pre_bl98_out pre_bl99_out
+ pre_bl100_out pre_bl101_out pre_bl102_out pre_bl103_out pre_bl104_out
+ pre_bl105_out pre_bl106_out pre_bl107_out pre_bl108_out pre_bl109_out
+ pre_bl110_out pre_bl111_out pre_bl112_out pre_bl113_out pre_bl114_out
+ pre_bl115_out pre_bl116_out pre_bl117_out pre_bl118_out pre_bl119_out
+ pre_bl120_out pre_bl121_out pre_bl122_out pre_bl123_out pre_bl124_out
+ pre_bl125_out pre_bl126_out pre_bl127_out pre_bl128_out pre_bl129_out
+ pre_bl130_out pre_bl131_out pre_bl132_out pre_bl133_out pre_bl134_out
+ pre_bl135_out pre_bl136_out pre_bl137_out pre_bl138_out pre_bl139_out
+ pre_bl140_out pre_bl141_out pre_bl142_out pre_bl143_out pre_bl144_out
+ pre_bl145_out pre_bl146_out pre_bl147_out pre_bl148_out pre_bl149_out
+ pre_bl150_out pre_bl151_out pre_bl152_out pre_bl153_out pre_bl154_out
+ pre_bl155_out pre_bl156_out pre_bl157_out pre_bl158_out pre_bl159_out
+ pre_bl160_out pre_bl161_out pre_bl162_out pre_bl163_out pre_bl164_out
+ pre_bl165_out pre_bl166_out pre_bl167_out pre_bl168_out pre_bl169_out
+ pre_bl170_out pre_bl171_out pre_bl172_out pre_bl173_out pre_bl174_out
+ pre_bl175_out pre_bl176_out pre_bl177_out pre_bl178_out pre_bl179_out
+ pre_bl180_out pre_bl181_out pre_bl182_out pre_bl183_out gate vdd
* OUTPUT: pre_bl0_out 
* OUTPUT: pre_bl1_out 
* OUTPUT: pre_bl2_out 
* OUTPUT: pre_bl3_out 
* OUTPUT: pre_bl4_out 
* OUTPUT: pre_bl5_out 
* OUTPUT: pre_bl6_out 
* OUTPUT: pre_bl7_out 
* OUTPUT: pre_bl8_out 
* OUTPUT: pre_bl9_out 
* OUTPUT: pre_bl10_out 
* OUTPUT: pre_bl11_out 
* OUTPUT: pre_bl12_out 
* OUTPUT: pre_bl13_out 
* OUTPUT: pre_bl14_out 
* OUTPUT: pre_bl15_out 
* OUTPUT: pre_bl16_out 
* OUTPUT: pre_bl17_out 
* OUTPUT: pre_bl18_out 
* OUTPUT: pre_bl19_out 
* OUTPUT: pre_bl20_out 
* OUTPUT: pre_bl21_out 
* OUTPUT: pre_bl22_out 
* OUTPUT: pre_bl23_out 
* OUTPUT: pre_bl24_out 
* OUTPUT: pre_bl25_out 
* OUTPUT: pre_bl26_out 
* OUTPUT: pre_bl27_out 
* OUTPUT: pre_bl28_out 
* OUTPUT: pre_bl29_out 
* OUTPUT: pre_bl30_out 
* OUTPUT: pre_bl31_out 
* OUTPUT: pre_bl32_out 
* OUTPUT: pre_bl33_out 
* OUTPUT: pre_bl34_out 
* OUTPUT: pre_bl35_out 
* OUTPUT: pre_bl36_out 
* OUTPUT: pre_bl37_out 
* OUTPUT: pre_bl38_out 
* OUTPUT: pre_bl39_out 
* OUTPUT: pre_bl40_out 
* OUTPUT: pre_bl41_out 
* OUTPUT: pre_bl42_out 
* OUTPUT: pre_bl43_out 
* OUTPUT: pre_bl44_out 
* OUTPUT: pre_bl45_out 
* OUTPUT: pre_bl46_out 
* OUTPUT: pre_bl47_out 
* OUTPUT: pre_bl48_out 
* OUTPUT: pre_bl49_out 
* OUTPUT: pre_bl50_out 
* OUTPUT: pre_bl51_out 
* OUTPUT: pre_bl52_out 
* OUTPUT: pre_bl53_out 
* OUTPUT: pre_bl54_out 
* OUTPUT: pre_bl55_out 
* OUTPUT: pre_bl56_out 
* OUTPUT: pre_bl57_out 
* OUTPUT: pre_bl58_out 
* OUTPUT: pre_bl59_out 
* OUTPUT: pre_bl60_out 
* OUTPUT: pre_bl61_out 
* OUTPUT: pre_bl62_out 
* OUTPUT: pre_bl63_out 
* OUTPUT: pre_bl64_out 
* OUTPUT: pre_bl65_out 
* OUTPUT: pre_bl66_out 
* OUTPUT: pre_bl67_out 
* OUTPUT: pre_bl68_out 
* OUTPUT: pre_bl69_out 
* OUTPUT: pre_bl70_out 
* OUTPUT: pre_bl71_out 
* OUTPUT: pre_bl72_out 
* OUTPUT: pre_bl73_out 
* OUTPUT: pre_bl74_out 
* OUTPUT: pre_bl75_out 
* OUTPUT: pre_bl76_out 
* OUTPUT: pre_bl77_out 
* OUTPUT: pre_bl78_out 
* OUTPUT: pre_bl79_out 
* OUTPUT: pre_bl80_out 
* OUTPUT: pre_bl81_out 
* OUTPUT: pre_bl82_out 
* OUTPUT: pre_bl83_out 
* OUTPUT: pre_bl84_out 
* OUTPUT: pre_bl85_out 
* OUTPUT: pre_bl86_out 
* OUTPUT: pre_bl87_out 
* OUTPUT: pre_bl88_out 
* OUTPUT: pre_bl89_out 
* OUTPUT: pre_bl90_out 
* OUTPUT: pre_bl91_out 
* OUTPUT: pre_bl92_out 
* OUTPUT: pre_bl93_out 
* OUTPUT: pre_bl94_out 
* OUTPUT: pre_bl95_out 
* OUTPUT: pre_bl96_out 
* OUTPUT: pre_bl97_out 
* OUTPUT: pre_bl98_out 
* OUTPUT: pre_bl99_out 
* OUTPUT: pre_bl100_out 
* OUTPUT: pre_bl101_out 
* OUTPUT: pre_bl102_out 
* OUTPUT: pre_bl103_out 
* OUTPUT: pre_bl104_out 
* OUTPUT: pre_bl105_out 
* OUTPUT: pre_bl106_out 
* OUTPUT: pre_bl107_out 
* OUTPUT: pre_bl108_out 
* OUTPUT: pre_bl109_out 
* OUTPUT: pre_bl110_out 
* OUTPUT: pre_bl111_out 
* OUTPUT: pre_bl112_out 
* OUTPUT: pre_bl113_out 
* OUTPUT: pre_bl114_out 
* OUTPUT: pre_bl115_out 
* OUTPUT: pre_bl116_out 
* OUTPUT: pre_bl117_out 
* OUTPUT: pre_bl118_out 
* OUTPUT: pre_bl119_out 
* OUTPUT: pre_bl120_out 
* OUTPUT: pre_bl121_out 
* OUTPUT: pre_bl122_out 
* OUTPUT: pre_bl123_out 
* OUTPUT: pre_bl124_out 
* OUTPUT: pre_bl125_out 
* OUTPUT: pre_bl126_out 
* OUTPUT: pre_bl127_out 
* OUTPUT: pre_bl128_out 
* OUTPUT: pre_bl129_out 
* OUTPUT: pre_bl130_out 
* OUTPUT: pre_bl131_out 
* OUTPUT: pre_bl132_out 
* OUTPUT: pre_bl133_out 
* OUTPUT: pre_bl134_out 
* OUTPUT: pre_bl135_out 
* OUTPUT: pre_bl136_out 
* OUTPUT: pre_bl137_out 
* OUTPUT: pre_bl138_out 
* OUTPUT: pre_bl139_out 
* OUTPUT: pre_bl140_out 
* OUTPUT: pre_bl141_out 
* OUTPUT: pre_bl142_out 
* OUTPUT: pre_bl143_out 
* OUTPUT: pre_bl144_out 
* OUTPUT: pre_bl145_out 
* OUTPUT: pre_bl146_out 
* OUTPUT: pre_bl147_out 
* OUTPUT: pre_bl148_out 
* OUTPUT: pre_bl149_out 
* OUTPUT: pre_bl150_out 
* OUTPUT: pre_bl151_out 
* OUTPUT: pre_bl152_out 
* OUTPUT: pre_bl153_out 
* OUTPUT: pre_bl154_out 
* OUTPUT: pre_bl155_out 
* OUTPUT: pre_bl156_out 
* OUTPUT: pre_bl157_out 
* OUTPUT: pre_bl158_out 
* OUTPUT: pre_bl159_out 
* OUTPUT: pre_bl160_out 
* OUTPUT: pre_bl161_out 
* OUTPUT: pre_bl162_out 
* OUTPUT: pre_bl163_out 
* OUTPUT: pre_bl164_out 
* OUTPUT: pre_bl165_out 
* OUTPUT: pre_bl166_out 
* OUTPUT: pre_bl167_out 
* OUTPUT: pre_bl168_out 
* OUTPUT: pre_bl169_out 
* OUTPUT: pre_bl170_out 
* OUTPUT: pre_bl171_out 
* OUTPUT: pre_bl172_out 
* OUTPUT: pre_bl173_out 
* OUTPUT: pre_bl174_out 
* OUTPUT: pre_bl175_out 
* OUTPUT: pre_bl176_out 
* OUTPUT: pre_bl177_out 
* OUTPUT: pre_bl178_out 
* OUTPUT: pre_bl179_out 
* OUTPUT: pre_bl180_out 
* OUTPUT: pre_bl181_out 
* OUTPUT: pre_bl182_out 
* OUTPUT: pre_bl183_out 
* INPUT : gate 
* POWER : vdd 
Xpmos_c0
+ vdd gate pre_bl0_out
+ sram_precharge_cell
Xpmos_c1
+ vdd gate pre_bl1_out
+ sram_precharge_cell
Xpmos_c2
+ vdd gate pre_bl2_out
+ sram_precharge_cell
Xpmos_c3
+ vdd gate pre_bl3_out
+ sram_precharge_cell
Xpmos_c4
+ vdd gate pre_bl4_out
+ sram_precharge_cell
Xpmos_c5
+ vdd gate pre_bl5_out
+ sram_precharge_cell
Xpmos_c6
+ vdd gate pre_bl6_out
+ sram_precharge_cell
Xpmos_c7
+ vdd gate pre_bl7_out
+ sram_precharge_cell
Xpmos_c8
+ vdd gate pre_bl8_out
+ sram_precharge_cell
Xpmos_c9
+ vdd gate pre_bl9_out
+ sram_precharge_cell
Xpmos_c10
+ vdd gate pre_bl10_out
+ sram_precharge_cell
Xpmos_c11
+ vdd gate pre_bl11_out
+ sram_precharge_cell
Xpmos_c12
+ vdd gate pre_bl12_out
+ sram_precharge_cell
Xpmos_c13
+ vdd gate pre_bl13_out
+ sram_precharge_cell
Xpmos_c14
+ vdd gate pre_bl14_out
+ sram_precharge_cell
Xpmos_c15
+ vdd gate pre_bl15_out
+ sram_precharge_cell
Xpmos_c16
+ vdd gate pre_bl16_out
+ sram_precharge_cell
Xpmos_c17
+ vdd gate pre_bl17_out
+ sram_precharge_cell
Xpmos_c18
+ vdd gate pre_bl18_out
+ sram_precharge_cell
Xpmos_c19
+ vdd gate pre_bl19_out
+ sram_precharge_cell
Xpmos_c20
+ vdd gate pre_bl20_out
+ sram_precharge_cell
Xpmos_c21
+ vdd gate pre_bl21_out
+ sram_precharge_cell
Xpmos_c22
+ vdd gate pre_bl22_out
+ sram_precharge_cell
Xpmos_c23
+ vdd gate pre_bl23_out
+ sram_precharge_cell
Xpmos_c24
+ vdd gate pre_bl24_out
+ sram_precharge_cell
Xpmos_c25
+ vdd gate pre_bl25_out
+ sram_precharge_cell
Xpmos_c26
+ vdd gate pre_bl26_out
+ sram_precharge_cell
Xpmos_c27
+ vdd gate pre_bl27_out
+ sram_precharge_cell
Xpmos_c28
+ vdd gate pre_bl28_out
+ sram_precharge_cell
Xpmos_c29
+ vdd gate pre_bl29_out
+ sram_precharge_cell
Xpmos_c30
+ vdd gate pre_bl30_out
+ sram_precharge_cell
Xpmos_c31
+ vdd gate pre_bl31_out
+ sram_precharge_cell
Xpmos_c32
+ vdd gate pre_bl32_out
+ sram_precharge_cell
Xpmos_c33
+ vdd gate pre_bl33_out
+ sram_precharge_cell
Xpmos_c34
+ vdd gate pre_bl34_out
+ sram_precharge_cell
Xpmos_c35
+ vdd gate pre_bl35_out
+ sram_precharge_cell
Xpmos_c36
+ vdd gate pre_bl36_out
+ sram_precharge_cell
Xpmos_c37
+ vdd gate pre_bl37_out
+ sram_precharge_cell
Xpmos_c38
+ vdd gate pre_bl38_out
+ sram_precharge_cell
Xpmos_c39
+ vdd gate pre_bl39_out
+ sram_precharge_cell
Xpmos_c40
+ vdd gate pre_bl40_out
+ sram_precharge_cell
Xpmos_c41
+ vdd gate pre_bl41_out
+ sram_precharge_cell
Xpmos_c42
+ vdd gate pre_bl42_out
+ sram_precharge_cell
Xpmos_c43
+ vdd gate pre_bl43_out
+ sram_precharge_cell
Xpmos_c44
+ vdd gate pre_bl44_out
+ sram_precharge_cell
Xpmos_c45
+ vdd gate pre_bl45_out
+ sram_precharge_cell
Xpmos_c46
+ vdd gate pre_bl46_out
+ sram_precharge_cell
Xpmos_c47
+ vdd gate pre_bl47_out
+ sram_precharge_cell
Xpmos_c48
+ vdd gate pre_bl48_out
+ sram_precharge_cell
Xpmos_c49
+ vdd gate pre_bl49_out
+ sram_precharge_cell
Xpmos_c50
+ vdd gate pre_bl50_out
+ sram_precharge_cell
Xpmos_c51
+ vdd gate pre_bl51_out
+ sram_precharge_cell
Xpmos_c52
+ vdd gate pre_bl52_out
+ sram_precharge_cell
Xpmos_c53
+ vdd gate pre_bl53_out
+ sram_precharge_cell
Xpmos_c54
+ vdd gate pre_bl54_out
+ sram_precharge_cell
Xpmos_c55
+ vdd gate pre_bl55_out
+ sram_precharge_cell
Xpmos_c56
+ vdd gate pre_bl56_out
+ sram_precharge_cell
Xpmos_c57
+ vdd gate pre_bl57_out
+ sram_precharge_cell
Xpmos_c58
+ vdd gate pre_bl58_out
+ sram_precharge_cell
Xpmos_c59
+ vdd gate pre_bl59_out
+ sram_precharge_cell
Xpmos_c60
+ vdd gate pre_bl60_out
+ sram_precharge_cell
Xpmos_c61
+ vdd gate pre_bl61_out
+ sram_precharge_cell
Xpmos_c62
+ vdd gate pre_bl62_out
+ sram_precharge_cell
Xpmos_c63
+ vdd gate pre_bl63_out
+ sram_precharge_cell
Xpmos_c64
+ vdd gate pre_bl64_out
+ sram_precharge_cell
Xpmos_c65
+ vdd gate pre_bl65_out
+ sram_precharge_cell
Xpmos_c66
+ vdd gate pre_bl66_out
+ sram_precharge_cell
Xpmos_c67
+ vdd gate pre_bl67_out
+ sram_precharge_cell
Xpmos_c68
+ vdd gate pre_bl68_out
+ sram_precharge_cell
Xpmos_c69
+ vdd gate pre_bl69_out
+ sram_precharge_cell
Xpmos_c70
+ vdd gate pre_bl70_out
+ sram_precharge_cell
Xpmos_c71
+ vdd gate pre_bl71_out
+ sram_precharge_cell
Xpmos_c72
+ vdd gate pre_bl72_out
+ sram_precharge_cell
Xpmos_c73
+ vdd gate pre_bl73_out
+ sram_precharge_cell
Xpmos_c74
+ vdd gate pre_bl74_out
+ sram_precharge_cell
Xpmos_c75
+ vdd gate pre_bl75_out
+ sram_precharge_cell
Xpmos_c76
+ vdd gate pre_bl76_out
+ sram_precharge_cell
Xpmos_c77
+ vdd gate pre_bl77_out
+ sram_precharge_cell
Xpmos_c78
+ vdd gate pre_bl78_out
+ sram_precharge_cell
Xpmos_c79
+ vdd gate pre_bl79_out
+ sram_precharge_cell
Xpmos_c80
+ vdd gate pre_bl80_out
+ sram_precharge_cell
Xpmos_c81
+ vdd gate pre_bl81_out
+ sram_precharge_cell
Xpmos_c82
+ vdd gate pre_bl82_out
+ sram_precharge_cell
Xpmos_c83
+ vdd gate pre_bl83_out
+ sram_precharge_cell
Xpmos_c84
+ vdd gate pre_bl84_out
+ sram_precharge_cell
Xpmos_c85
+ vdd gate pre_bl85_out
+ sram_precharge_cell
Xpmos_c86
+ vdd gate pre_bl86_out
+ sram_precharge_cell
Xpmos_c87
+ vdd gate pre_bl87_out
+ sram_precharge_cell
Xpmos_c88
+ vdd gate pre_bl88_out
+ sram_precharge_cell
Xpmos_c89
+ vdd gate pre_bl89_out
+ sram_precharge_cell
Xpmos_c90
+ vdd gate pre_bl90_out
+ sram_precharge_cell
Xpmos_c91
+ vdd gate pre_bl91_out
+ sram_precharge_cell
Xpmos_c92
+ vdd gate pre_bl92_out
+ sram_precharge_cell
Xpmos_c93
+ vdd gate pre_bl93_out
+ sram_precharge_cell
Xpmos_c94
+ vdd gate pre_bl94_out
+ sram_precharge_cell
Xpmos_c95
+ vdd gate pre_bl95_out
+ sram_precharge_cell
Xpmos_c96
+ vdd gate pre_bl96_out
+ sram_precharge_cell
Xpmos_c97
+ vdd gate pre_bl97_out
+ sram_precharge_cell
Xpmos_c98
+ vdd gate pre_bl98_out
+ sram_precharge_cell
Xpmos_c99
+ vdd gate pre_bl99_out
+ sram_precharge_cell
Xpmos_c100
+ vdd gate pre_bl100_out
+ sram_precharge_cell
Xpmos_c101
+ vdd gate pre_bl101_out
+ sram_precharge_cell
Xpmos_c102
+ vdd gate pre_bl102_out
+ sram_precharge_cell
Xpmos_c103
+ vdd gate pre_bl103_out
+ sram_precharge_cell
Xpmos_c104
+ vdd gate pre_bl104_out
+ sram_precharge_cell
Xpmos_c105
+ vdd gate pre_bl105_out
+ sram_precharge_cell
Xpmos_c106
+ vdd gate pre_bl106_out
+ sram_precharge_cell
Xpmos_c107
+ vdd gate pre_bl107_out
+ sram_precharge_cell
Xpmos_c108
+ vdd gate pre_bl108_out
+ sram_precharge_cell
Xpmos_c109
+ vdd gate pre_bl109_out
+ sram_precharge_cell
Xpmos_c110
+ vdd gate pre_bl110_out
+ sram_precharge_cell
Xpmos_c111
+ vdd gate pre_bl111_out
+ sram_precharge_cell
Xpmos_c112
+ vdd gate pre_bl112_out
+ sram_precharge_cell
Xpmos_c113
+ vdd gate pre_bl113_out
+ sram_precharge_cell
Xpmos_c114
+ vdd gate pre_bl114_out
+ sram_precharge_cell
Xpmos_c115
+ vdd gate pre_bl115_out
+ sram_precharge_cell
Xpmos_c116
+ vdd gate pre_bl116_out
+ sram_precharge_cell
Xpmos_c117
+ vdd gate pre_bl117_out
+ sram_precharge_cell
Xpmos_c118
+ vdd gate pre_bl118_out
+ sram_precharge_cell
Xpmos_c119
+ vdd gate pre_bl119_out
+ sram_precharge_cell
Xpmos_c120
+ vdd gate pre_bl120_out
+ sram_precharge_cell
Xpmos_c121
+ vdd gate pre_bl121_out
+ sram_precharge_cell
Xpmos_c122
+ vdd gate pre_bl122_out
+ sram_precharge_cell
Xpmos_c123
+ vdd gate pre_bl123_out
+ sram_precharge_cell
Xpmos_c124
+ vdd gate pre_bl124_out
+ sram_precharge_cell
Xpmos_c125
+ vdd gate pre_bl125_out
+ sram_precharge_cell
Xpmos_c126
+ vdd gate pre_bl126_out
+ sram_precharge_cell
Xpmos_c127
+ vdd gate pre_bl127_out
+ sram_precharge_cell
Xpmos_c128
+ vdd gate pre_bl128_out
+ sram_precharge_cell
Xpmos_c129
+ vdd gate pre_bl129_out
+ sram_precharge_cell
Xpmos_c130
+ vdd gate pre_bl130_out
+ sram_precharge_cell
Xpmos_c131
+ vdd gate pre_bl131_out
+ sram_precharge_cell
Xpmos_c132
+ vdd gate pre_bl132_out
+ sram_precharge_cell
Xpmos_c133
+ vdd gate pre_bl133_out
+ sram_precharge_cell
Xpmos_c134
+ vdd gate pre_bl134_out
+ sram_precharge_cell
Xpmos_c135
+ vdd gate pre_bl135_out
+ sram_precharge_cell
Xpmos_c136
+ vdd gate pre_bl136_out
+ sram_precharge_cell
Xpmos_c137
+ vdd gate pre_bl137_out
+ sram_precharge_cell
Xpmos_c138
+ vdd gate pre_bl138_out
+ sram_precharge_cell
Xpmos_c139
+ vdd gate pre_bl139_out
+ sram_precharge_cell
Xpmos_c140
+ vdd gate pre_bl140_out
+ sram_precharge_cell
Xpmos_c141
+ vdd gate pre_bl141_out
+ sram_precharge_cell
Xpmos_c142
+ vdd gate pre_bl142_out
+ sram_precharge_cell
Xpmos_c143
+ vdd gate pre_bl143_out
+ sram_precharge_cell
Xpmos_c144
+ vdd gate pre_bl144_out
+ sram_precharge_cell
Xpmos_c145
+ vdd gate pre_bl145_out
+ sram_precharge_cell
Xpmos_c146
+ vdd gate pre_bl146_out
+ sram_precharge_cell
Xpmos_c147
+ vdd gate pre_bl147_out
+ sram_precharge_cell
Xpmos_c148
+ vdd gate pre_bl148_out
+ sram_precharge_cell
Xpmos_c149
+ vdd gate pre_bl149_out
+ sram_precharge_cell
Xpmos_c150
+ vdd gate pre_bl150_out
+ sram_precharge_cell
Xpmos_c151
+ vdd gate pre_bl151_out
+ sram_precharge_cell
Xpmos_c152
+ vdd gate pre_bl152_out
+ sram_precharge_cell
Xpmos_c153
+ vdd gate pre_bl153_out
+ sram_precharge_cell
Xpmos_c154
+ vdd gate pre_bl154_out
+ sram_precharge_cell
Xpmos_c155
+ vdd gate pre_bl155_out
+ sram_precharge_cell
Xpmos_c156
+ vdd gate pre_bl156_out
+ sram_precharge_cell
Xpmos_c157
+ vdd gate pre_bl157_out
+ sram_precharge_cell
Xpmos_c158
+ vdd gate pre_bl158_out
+ sram_precharge_cell
Xpmos_c159
+ vdd gate pre_bl159_out
+ sram_precharge_cell
Xpmos_c160
+ vdd gate pre_bl160_out
+ sram_precharge_cell
Xpmos_c161
+ vdd gate pre_bl161_out
+ sram_precharge_cell
Xpmos_c162
+ vdd gate pre_bl162_out
+ sram_precharge_cell
Xpmos_c163
+ vdd gate pre_bl163_out
+ sram_precharge_cell
Xpmos_c164
+ vdd gate pre_bl164_out
+ sram_precharge_cell
Xpmos_c165
+ vdd gate pre_bl165_out
+ sram_precharge_cell
Xpmos_c166
+ vdd gate pre_bl166_out
+ sram_precharge_cell
Xpmos_c167
+ vdd gate pre_bl167_out
+ sram_precharge_cell
Xpmos_c168
+ vdd gate pre_bl168_out
+ sram_precharge_cell
Xpmos_c169
+ vdd gate pre_bl169_out
+ sram_precharge_cell
Xpmos_c170
+ vdd gate pre_bl170_out
+ sram_precharge_cell
Xpmos_c171
+ vdd gate pre_bl171_out
+ sram_precharge_cell
Xpmos_c172
+ vdd gate pre_bl172_out
+ sram_precharge_cell
Xpmos_c173
+ vdd gate pre_bl173_out
+ sram_precharge_cell
Xpmos_c174
+ vdd gate pre_bl174_out
+ sram_precharge_cell
Xpmos_c175
+ vdd gate pre_bl175_out
+ sram_precharge_cell
Xpmos_c176
+ vdd gate pre_bl176_out
+ sram_precharge_cell
Xpmos_c177
+ vdd gate pre_bl177_out
+ sram_precharge_cell
Xpmos_c178
+ vdd gate pre_bl178_out
+ sram_precharge_cell
Xpmos_c179
+ vdd gate pre_bl179_out
+ sram_precharge_cell
Xpmos_c180
+ vdd gate pre_bl180_out
+ sram_precharge_cell
Xpmos_c181
+ vdd gate pre_bl181_out
+ sram_precharge_cell
Xpmos_c182
+ vdd gate pre_bl182_out
+ sram_precharge_cell
Xpmos_c183
+ vdd gate pre_bl183_out
+ sram_precharge_cell
.ENDS sram_rom_precharge_array

.SUBCKT sram_rom_base_array
+ bl_0_0 bl_0_1 bl_0_2 bl_0_3 bl_0_4 bl_0_5 bl_0_6 bl_0_7 bl_0_8 bl_0_9
+ bl_0_10 bl_0_11 bl_0_12 bl_0_13 bl_0_14 bl_0_15 bl_0_16 bl_0_17
+ bl_0_18 bl_0_19 bl_0_20 bl_0_21 bl_0_22 bl_0_23 bl_0_24 bl_0_25
+ bl_0_26 bl_0_27 bl_0_28 bl_0_29 bl_0_30 bl_0_31 bl_0_32 bl_0_33
+ bl_0_34 bl_0_35 bl_0_36 bl_0_37 bl_0_38 bl_0_39 bl_0_40 bl_0_41
+ bl_0_42 bl_0_43 bl_0_44 bl_0_45 bl_0_46 bl_0_47 bl_0_48 bl_0_49
+ bl_0_50 bl_0_51 bl_0_52 bl_0_53 bl_0_54 bl_0_55 bl_0_56 bl_0_57
+ bl_0_58 bl_0_59 bl_0_60 bl_0_61 bl_0_62 bl_0_63 bl_0_64 bl_0_65
+ bl_0_66 bl_0_67 bl_0_68 bl_0_69 bl_0_70 bl_0_71 bl_0_72 bl_0_73
+ bl_0_74 bl_0_75 bl_0_76 bl_0_77 bl_0_78 bl_0_79 bl_0_80 bl_0_81
+ bl_0_82 bl_0_83 bl_0_84 bl_0_85 bl_0_86 bl_0_87 bl_0_88 bl_0_89
+ bl_0_90 bl_0_91 bl_0_92 bl_0_93 bl_0_94 bl_0_95 bl_0_96 bl_0_97
+ bl_0_98 bl_0_99 bl_0_100 bl_0_101 bl_0_102 bl_0_103 bl_0_104 bl_0_105
+ bl_0_106 bl_0_107 bl_0_108 bl_0_109 bl_0_110 bl_0_111 bl_0_112
+ bl_0_113 bl_0_114 bl_0_115 bl_0_116 bl_0_117 bl_0_118 bl_0_119
+ bl_0_120 bl_0_121 bl_0_122 bl_0_123 bl_0_124 bl_0_125 bl_0_126
+ bl_0_127 bl_0_128 bl_0_129 bl_0_130 bl_0_131 bl_0_132 bl_0_133
+ bl_0_134 bl_0_135 bl_0_136 bl_0_137 bl_0_138 bl_0_139 bl_0_140
+ bl_0_141 bl_0_142 bl_0_143 bl_0_144 bl_0_145 bl_0_146 bl_0_147
+ bl_0_148 bl_0_149 bl_0_150 bl_0_151 bl_0_152 bl_0_153 bl_0_154
+ bl_0_155 bl_0_156 bl_0_157 bl_0_158 bl_0_159 bl_0_160 bl_0_161
+ bl_0_162 bl_0_163 bl_0_164 bl_0_165 bl_0_166 bl_0_167 bl_0_168
+ bl_0_169 bl_0_170 bl_0_171 bl_0_172 bl_0_173 bl_0_174 bl_0_175
+ bl_0_176 bl_0_177 bl_0_178 bl_0_179 bl_0_180 bl_0_181 bl_0_182
+ bl_0_183 wl_0_0 wl_0_1 wl_0_2 wl_0_3 wl_0_4 wl_0_5 wl_0_6 wl_0_7
+ wl_0_8 wl_0_9 wl_0_10 wl_0_11 wl_0_12 wl_0_13 wl_0_14 wl_0_15 wl_0_16
+ wl_0_17 wl_0_18 wl_0_19 wl_0_20 wl_0_21 wl_0_22 wl_0_23 wl_0_24
+ wl_0_25 wl_0_26 wl_0_27 wl_0_28 wl_0_29 wl_0_30 wl_0_31 wl_0_32
+ wl_0_33 wl_0_34 wl_0_35 wl_0_36 wl_0_37 wl_0_38 wl_0_39 wl_0_40
+ wl_0_41 wl_0_42 wl_0_43 wl_0_44 wl_0_45 wl_0_46 wl_0_47 wl_0_48
+ wl_0_49 wl_0_50 wl_0_51 wl_0_52 wl_0_53 wl_0_54 wl_0_55 wl_0_56
+ wl_0_57 wl_0_58 wl_0_59 wl_0_60 wl_0_61 wl_0_62 wl_0_63 wl_0_64
+ wl_0_65 wl_0_66 wl_0_67 wl_0_68 wl_0_69 wl_0_70 wl_0_71 wl_0_72
+ wl_0_73 wl_0_74 wl_0_75 wl_0_76 wl_0_77 wl_0_78 wl_0_79 wl_0_80
+ wl_0_81 wl_0_82 wl_0_83 wl_0_84 wl_0_85 wl_0_86 wl_0_87 wl_0_88
+ precharge vdd gnd
* OUTPUT: bl_0_0 
* OUTPUT: bl_0_1 
* OUTPUT: bl_0_2 
* OUTPUT: bl_0_3 
* OUTPUT: bl_0_4 
* OUTPUT: bl_0_5 
* OUTPUT: bl_0_6 
* OUTPUT: bl_0_7 
* OUTPUT: bl_0_8 
* OUTPUT: bl_0_9 
* OUTPUT: bl_0_10 
* OUTPUT: bl_0_11 
* OUTPUT: bl_0_12 
* OUTPUT: bl_0_13 
* OUTPUT: bl_0_14 
* OUTPUT: bl_0_15 
* OUTPUT: bl_0_16 
* OUTPUT: bl_0_17 
* OUTPUT: bl_0_18 
* OUTPUT: bl_0_19 
* OUTPUT: bl_0_20 
* OUTPUT: bl_0_21 
* OUTPUT: bl_0_22 
* OUTPUT: bl_0_23 
* OUTPUT: bl_0_24 
* OUTPUT: bl_0_25 
* OUTPUT: bl_0_26 
* OUTPUT: bl_0_27 
* OUTPUT: bl_0_28 
* OUTPUT: bl_0_29 
* OUTPUT: bl_0_30 
* OUTPUT: bl_0_31 
* OUTPUT: bl_0_32 
* OUTPUT: bl_0_33 
* OUTPUT: bl_0_34 
* OUTPUT: bl_0_35 
* OUTPUT: bl_0_36 
* OUTPUT: bl_0_37 
* OUTPUT: bl_0_38 
* OUTPUT: bl_0_39 
* OUTPUT: bl_0_40 
* OUTPUT: bl_0_41 
* OUTPUT: bl_0_42 
* OUTPUT: bl_0_43 
* OUTPUT: bl_0_44 
* OUTPUT: bl_0_45 
* OUTPUT: bl_0_46 
* OUTPUT: bl_0_47 
* OUTPUT: bl_0_48 
* OUTPUT: bl_0_49 
* OUTPUT: bl_0_50 
* OUTPUT: bl_0_51 
* OUTPUT: bl_0_52 
* OUTPUT: bl_0_53 
* OUTPUT: bl_0_54 
* OUTPUT: bl_0_55 
* OUTPUT: bl_0_56 
* OUTPUT: bl_0_57 
* OUTPUT: bl_0_58 
* OUTPUT: bl_0_59 
* OUTPUT: bl_0_60 
* OUTPUT: bl_0_61 
* OUTPUT: bl_0_62 
* OUTPUT: bl_0_63 
* OUTPUT: bl_0_64 
* OUTPUT: bl_0_65 
* OUTPUT: bl_0_66 
* OUTPUT: bl_0_67 
* OUTPUT: bl_0_68 
* OUTPUT: bl_0_69 
* OUTPUT: bl_0_70 
* OUTPUT: bl_0_71 
* OUTPUT: bl_0_72 
* OUTPUT: bl_0_73 
* OUTPUT: bl_0_74 
* OUTPUT: bl_0_75 
* OUTPUT: bl_0_76 
* OUTPUT: bl_0_77 
* OUTPUT: bl_0_78 
* OUTPUT: bl_0_79 
* OUTPUT: bl_0_80 
* OUTPUT: bl_0_81 
* OUTPUT: bl_0_82 
* OUTPUT: bl_0_83 
* OUTPUT: bl_0_84 
* OUTPUT: bl_0_85 
* OUTPUT: bl_0_86 
* OUTPUT: bl_0_87 
* OUTPUT: bl_0_88 
* OUTPUT: bl_0_89 
* OUTPUT: bl_0_90 
* OUTPUT: bl_0_91 
* OUTPUT: bl_0_92 
* OUTPUT: bl_0_93 
* OUTPUT: bl_0_94 
* OUTPUT: bl_0_95 
* OUTPUT: bl_0_96 
* OUTPUT: bl_0_97 
* OUTPUT: bl_0_98 
* OUTPUT: bl_0_99 
* OUTPUT: bl_0_100 
* OUTPUT: bl_0_101 
* OUTPUT: bl_0_102 
* OUTPUT: bl_0_103 
* OUTPUT: bl_0_104 
* OUTPUT: bl_0_105 
* OUTPUT: bl_0_106 
* OUTPUT: bl_0_107 
* OUTPUT: bl_0_108 
* OUTPUT: bl_0_109 
* OUTPUT: bl_0_110 
* OUTPUT: bl_0_111 
* OUTPUT: bl_0_112 
* OUTPUT: bl_0_113 
* OUTPUT: bl_0_114 
* OUTPUT: bl_0_115 
* OUTPUT: bl_0_116 
* OUTPUT: bl_0_117 
* OUTPUT: bl_0_118 
* OUTPUT: bl_0_119 
* OUTPUT: bl_0_120 
* OUTPUT: bl_0_121 
* OUTPUT: bl_0_122 
* OUTPUT: bl_0_123 
* OUTPUT: bl_0_124 
* OUTPUT: bl_0_125 
* OUTPUT: bl_0_126 
* OUTPUT: bl_0_127 
* OUTPUT: bl_0_128 
* OUTPUT: bl_0_129 
* OUTPUT: bl_0_130 
* OUTPUT: bl_0_131 
* OUTPUT: bl_0_132 
* OUTPUT: bl_0_133 
* OUTPUT: bl_0_134 
* OUTPUT: bl_0_135 
* OUTPUT: bl_0_136 
* OUTPUT: bl_0_137 
* OUTPUT: bl_0_138 
* OUTPUT: bl_0_139 
* OUTPUT: bl_0_140 
* OUTPUT: bl_0_141 
* OUTPUT: bl_0_142 
* OUTPUT: bl_0_143 
* OUTPUT: bl_0_144 
* OUTPUT: bl_0_145 
* OUTPUT: bl_0_146 
* OUTPUT: bl_0_147 
* OUTPUT: bl_0_148 
* OUTPUT: bl_0_149 
* OUTPUT: bl_0_150 
* OUTPUT: bl_0_151 
* OUTPUT: bl_0_152 
* OUTPUT: bl_0_153 
* OUTPUT: bl_0_154 
* OUTPUT: bl_0_155 
* OUTPUT: bl_0_156 
* OUTPUT: bl_0_157 
* OUTPUT: bl_0_158 
* OUTPUT: bl_0_159 
* OUTPUT: bl_0_160 
* OUTPUT: bl_0_161 
* OUTPUT: bl_0_162 
* OUTPUT: bl_0_163 
* OUTPUT: bl_0_164 
* OUTPUT: bl_0_165 
* OUTPUT: bl_0_166 
* OUTPUT: bl_0_167 
* OUTPUT: bl_0_168 
* OUTPUT: bl_0_169 
* OUTPUT: bl_0_170 
* OUTPUT: bl_0_171 
* OUTPUT: bl_0_172 
* OUTPUT: bl_0_173 
* OUTPUT: bl_0_174 
* OUTPUT: bl_0_175 
* OUTPUT: bl_0_176 
* OUTPUT: bl_0_177 
* OUTPUT: bl_0_178 
* OUTPUT: bl_0_179 
* OUTPUT: bl_0_180 
* OUTPUT: bl_0_181 
* OUTPUT: bl_0_182 
* OUTPUT: bl_0_183 
* INPUT : wl_0_0 
* INPUT : wl_0_1 
* INPUT : wl_0_2 
* INPUT : wl_0_3 
* INPUT : wl_0_4 
* INPUT : wl_0_5 
* INPUT : wl_0_6 
* INPUT : wl_0_7 
* INPUT : wl_0_8 
* INPUT : wl_0_9 
* INPUT : wl_0_10 
* INPUT : wl_0_11 
* INPUT : wl_0_12 
* INPUT : wl_0_13 
* INPUT : wl_0_14 
* INPUT : wl_0_15 
* INPUT : wl_0_16 
* INPUT : wl_0_17 
* INPUT : wl_0_18 
* INPUT : wl_0_19 
* INPUT : wl_0_20 
* INPUT : wl_0_21 
* INPUT : wl_0_22 
* INPUT : wl_0_23 
* INPUT : wl_0_24 
* INPUT : wl_0_25 
* INPUT : wl_0_26 
* INPUT : wl_0_27 
* INPUT : wl_0_28 
* INPUT : wl_0_29 
* INPUT : wl_0_30 
* INPUT : wl_0_31 
* INPUT : wl_0_32 
* INPUT : wl_0_33 
* INPUT : wl_0_34 
* INPUT : wl_0_35 
* INPUT : wl_0_36 
* INPUT : wl_0_37 
* INPUT : wl_0_38 
* INPUT : wl_0_39 
* INPUT : wl_0_40 
* INPUT : wl_0_41 
* INPUT : wl_0_42 
* INPUT : wl_0_43 
* INPUT : wl_0_44 
* INPUT : wl_0_45 
* INPUT : wl_0_46 
* INPUT : wl_0_47 
* INPUT : wl_0_48 
* INPUT : wl_0_49 
* INPUT : wl_0_50 
* INPUT : wl_0_51 
* INPUT : wl_0_52 
* INPUT : wl_0_53 
* INPUT : wl_0_54 
* INPUT : wl_0_55 
* INPUT : wl_0_56 
* INPUT : wl_0_57 
* INPUT : wl_0_58 
* INPUT : wl_0_59 
* INPUT : wl_0_60 
* INPUT : wl_0_61 
* INPUT : wl_0_62 
* INPUT : wl_0_63 
* INPUT : wl_0_64 
* INPUT : wl_0_65 
* INPUT : wl_0_66 
* INPUT : wl_0_67 
* INPUT : wl_0_68 
* INPUT : wl_0_69 
* INPUT : wl_0_70 
* INPUT : wl_0_71 
* INPUT : wl_0_72 
* INPUT : wl_0_73 
* INPUT : wl_0_74 
* INPUT : wl_0_75 
* INPUT : wl_0_76 
* INPUT : wl_0_77 
* INPUT : wl_0_78 
* INPUT : wl_0_79 
* INPUT : wl_0_80 
* INPUT : wl_0_81 
* INPUT : wl_0_82 
* INPUT : wl_0_83 
* INPUT : wl_0_84 
* INPUT : wl_0_85 
* INPUT : wl_0_86 
* INPUT : wl_0_87 
* INPUT : wl_0_88 
* INPUT : precharge 
* POWER : vdd 
* GROUND: gnd 
Xbit_r0_c0
+ bl_int_0_0 bl_0_0 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c1
+ bl_int_0_1 bl_0_1 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c2
+ bl_int_0_2 bl_0_2 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c3
+ bl_int_0_3 bl_0_3 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c4
+ bl_int_0_4 bl_0_4 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c5
+ bl_int_0_5 bl_0_5 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c6
+ bl_int_0_6 bl_0_6 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c7
+ bl_int_0_7 bl_0_7 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c8
+ bl_int_0_8 bl_0_8 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c9
+ bl_int_0_9 bl_0_9 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c10
+ bl_int_0_10 bl_0_10 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c11
+ bl_int_0_11 bl_0_11 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c12
+ bl_int_0_12 bl_0_12 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c13
+ bl_int_0_13 bl_0_13 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c14
+ bl_int_0_14 bl_0_14 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c15
+ bl_int_0_15 bl_0_15 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c16
+ bl_int_0_16 bl_0_16 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c17
+ bl_int_0_17 bl_0_17 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c18
+ bl_int_0_18 bl_0_18 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c19
+ bl_int_0_19 bl_0_19 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c20
+ bl_int_0_20 bl_0_20 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c21
+ bl_int_0_21 bl_0_21 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c22
+ bl_int_0_22 bl_0_22 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c23
+ bl_int_0_23 bl_0_23 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c24
+ bl_int_0_24 bl_0_24 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c25
+ bl_int_0_25 bl_0_25 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c26
+ bl_int_0_26 bl_0_26 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c27
+ bl_int_0_27 bl_0_27 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c28
+ bl_int_0_28 bl_0_28 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c29
+ bl_int_0_29 bl_0_29 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c30
+ bl_int_0_30 bl_0_30 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c31
+ bl_int_0_31 bl_0_31 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c32
+ bl_int_0_32 bl_0_32 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c33
+ bl_int_0_33 bl_0_33 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c34
+ bl_int_0_34 bl_0_34 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c35
+ bl_int_0_35 bl_0_35 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c36
+ bl_int_0_36 bl_0_36 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c37
+ bl_int_0_37 bl_0_37 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c38
+ bl_int_0_38 bl_0_38 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c39
+ bl_int_0_39 bl_0_39 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c40
+ bl_int_0_40 bl_0_40 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c41
+ bl_int_0_41 bl_0_41 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c42
+ bl_int_0_42 bl_0_42 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c43
+ bl_int_0_43 bl_0_43 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c44
+ bl_int_0_44 bl_0_44 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c45
+ bl_int_0_45 bl_0_45 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c46
+ bl_int_0_46 bl_0_46 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c47
+ bl_int_0_47 bl_0_47 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c48
+ bl_int_0_48 bl_0_48 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c49
+ bl_int_0_49 bl_0_49 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c50
+ bl_int_0_50 bl_0_50 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c51
+ bl_int_0_51 bl_0_51 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c52
+ bl_int_0_52 bl_0_52 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c53
+ bl_int_0_53 bl_0_53 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c54
+ bl_int_0_54 bl_0_54 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c55
+ bl_int_0_55 bl_0_55 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c56
+ bl_int_0_56 bl_0_56 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c57
+ bl_int_0_57 bl_0_57 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c58
+ bl_int_0_58 bl_0_58 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c59
+ bl_int_0_59 bl_0_59 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c60
+ bl_int_0_60 bl_0_60 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c61
+ bl_int_0_61 bl_0_61 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c62
+ bl_int_0_62 bl_0_62 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c63
+ bl_int_0_63 bl_0_63 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c64
+ bl_int_0_64 bl_0_64 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c65
+ bl_int_0_65 bl_0_65 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c66
+ bl_int_0_66 bl_0_66 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c67
+ bl_int_0_67 bl_0_67 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c68
+ bl_int_0_68 bl_0_68 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c69
+ bl_int_0_69 bl_0_69 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c70
+ bl_int_0_70 bl_0_70 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c71
+ bl_int_0_71 bl_0_71 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c72
+ bl_int_0_72 bl_0_72 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c73
+ bl_int_0_73 bl_0_73 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c74
+ bl_int_0_74 bl_0_74 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c75
+ bl_int_0_75 bl_0_75 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c76
+ bl_int_0_76 bl_0_76 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c77
+ bl_int_0_77 bl_0_77 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c78
+ bl_int_0_78 bl_0_78 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c79
+ bl_int_0_79 bl_0_79 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c80
+ bl_int_0_80 bl_0_80 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c81
+ bl_int_0_81 bl_0_81 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c82
+ bl_int_0_82 bl_0_82 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c83
+ bl_int_0_83 bl_0_83 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c84
+ bl_int_0_84 bl_0_84 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c85
+ bl_int_0_85 bl_0_85 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c86
+ bl_int_0_86 bl_0_86 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c87
+ bl_int_0_87 bl_0_87 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c88
+ bl_int_0_88 bl_0_88 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c89
+ bl_int_0_89 bl_0_89 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c90
+ bl_int_0_90 bl_0_90 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c91
+ bl_int_0_91 bl_0_91 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c92
+ bl_int_0_92 bl_0_92 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c93
+ bl_int_0_93 bl_0_93 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c94
+ bl_int_0_94 bl_0_94 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c95
+ bl_int_0_95 bl_0_95 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c96
+ bl_int_0_96 bl_0_96 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c97
+ bl_int_0_97 bl_0_97 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c98
+ bl_int_0_98 bl_0_98 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c99
+ bl_int_0_99 bl_0_99 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c100
+ bl_int_0_100 bl_0_100 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c101
+ bl_int_0_101 bl_0_101 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c102
+ bl_int_0_102 bl_0_102 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c103
+ bl_int_0_103 bl_0_103 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c104
+ bl_int_0_104 bl_0_104 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c105
+ bl_int_0_105 bl_0_105 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c106
+ bl_int_0_106 bl_0_106 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c107
+ bl_int_0_107 bl_0_107 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c108
+ bl_int_0_108 bl_0_108 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c109
+ bl_int_0_109 bl_0_109 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c110
+ bl_int_0_110 bl_0_110 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c111
+ bl_int_0_111 bl_0_111 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c112
+ bl_int_0_112 bl_0_112 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c113
+ bl_int_0_113 bl_0_113 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c114
+ bl_int_0_114 bl_0_114 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c115
+ bl_int_0_115 bl_0_115 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c116
+ bl_int_0_116 bl_0_116 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c117
+ bl_int_0_117 bl_0_117 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c118
+ bl_int_0_118 bl_0_118 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c119
+ bl_int_0_119 bl_0_119 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c120
+ bl_int_0_120 bl_0_120 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c121
+ bl_int_0_121 bl_0_121 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c122
+ bl_int_0_122 bl_0_122 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c123
+ bl_int_0_123 bl_0_123 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c124
+ bl_int_0_124 bl_0_124 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c125
+ bl_int_0_125 bl_0_125 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c126
+ bl_int_0_126 bl_0_126 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c127
+ bl_int_0_127 bl_0_127 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c128
+ bl_int_0_128 bl_0_128 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c129
+ bl_int_0_129 bl_0_129 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c130
+ bl_int_0_130 bl_0_130 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c131
+ bl_int_0_131 bl_0_131 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c132
+ bl_int_0_132 bl_0_132 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c133
+ bl_int_0_133 bl_0_133 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c134
+ bl_int_0_134 bl_0_134 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c135
+ bl_int_0_135 bl_0_135 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c136
+ bl_int_0_136 bl_0_136 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c137
+ bl_int_0_137 bl_0_137 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c138
+ bl_int_0_138 bl_0_138 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c139
+ bl_int_0_139 bl_0_139 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c140
+ bl_int_0_140 bl_0_140 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c141
+ bl_int_0_141 bl_0_141 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c142
+ bl_int_0_142 bl_0_142 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c143
+ bl_int_0_143 bl_0_143 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c144
+ bl_int_0_144 bl_0_144 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c145
+ bl_int_0_145 bl_0_145 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c146
+ bl_int_0_146 bl_0_146 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c147
+ bl_int_0_147 bl_0_147 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c148
+ bl_int_0_148 bl_0_148 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c149
+ bl_int_0_149 bl_0_149 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c150
+ bl_int_0_150 bl_0_150 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c151
+ bl_int_0_151 bl_0_151 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c152
+ bl_int_0_152 bl_0_152 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c153
+ bl_int_0_153 bl_0_153 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c154
+ bl_int_0_154 bl_0_154 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c155
+ bl_int_0_155 bl_0_155 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c156
+ bl_int_0_156 bl_0_156 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c157
+ bl_int_0_157 bl_0_157 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c158
+ bl_int_0_158 bl_0_158 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c159
+ bl_int_0_159 bl_0_159 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c160
+ bl_int_0_160 bl_0_160 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c161
+ bl_int_0_161 bl_0_161 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c162
+ bl_int_0_162 bl_0_162 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c163
+ bl_int_0_163 bl_0_163 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c164
+ bl_int_0_164 bl_0_164 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c165
+ bl_int_0_165 bl_0_165 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c166
+ bl_int_0_166 bl_0_166 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c167
+ bl_int_0_167 bl_0_167 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c168
+ bl_int_0_168 bl_0_168 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c169
+ bl_int_0_169 bl_0_169 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c170
+ bl_int_0_170 bl_0_170 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c171
+ bl_int_0_171 bl_0_171 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c172
+ bl_int_0_172 bl_0_172 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c173
+ bl_int_0_173 bl_0_173 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c174
+ bl_int_0_174 bl_0_174 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c175
+ bl_int_0_175 bl_0_175 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c176
+ bl_int_0_176 bl_0_176 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c177
+ bl_int_0_177 bl_0_177 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c178
+ bl_int_0_178 bl_0_178 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c179
+ bl_int_0_179 bl_0_179 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c180
+ bl_int_0_180 bl_0_180 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c181
+ bl_int_0_181 bl_0_181 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c182
+ bl_int_0_182 bl_0_182 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r0_c183
+ bl_int_0_183 bl_0_183 wl_0_0 gnd
+ sram_rom_base_one_cell
Xbit_r1_c0
+ bl_int_1_0 bl_int_0_0 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c1
+ bl_int_1_1 bl_int_0_1 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c2
+ bl_int_1_2 bl_int_0_2 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c3
+ bl_int_1_3 bl_int_0_3 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c4
+ bl_int_1_4 bl_int_0_4 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c5
+ bl_int_1_5 bl_int_0_5 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c6
+ bl_int_1_6 bl_int_0_6 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c7
+ bl_int_1_7 bl_int_0_7 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c8
+ bl_int_1_8 bl_int_0_8 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c9
+ bl_int_1_9 bl_int_0_9 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c10
+ bl_int_1_10 bl_int_0_10 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c11
+ bl_int_1_11 bl_int_0_11 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c12
+ bl_int_1_12 bl_int_0_12 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c13
+ bl_int_1_13 bl_int_0_13 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c14
+ bl_int_1_14 bl_int_0_14 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c15
+ bl_int_1_15 bl_int_0_15 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c16
+ bl_int_1_16 bl_int_0_16 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c17
+ bl_int_1_17 bl_int_0_17 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c18
+ bl_int_1_18 bl_int_0_18 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c19
+ bl_int_1_19 bl_int_0_19 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c20
+ bl_int_1_20 bl_int_0_20 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c21
+ bl_int_1_21 bl_int_0_21 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c22
+ bl_int_1_22 bl_int_0_22 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c23
+ bl_int_1_23 bl_int_0_23 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c24
+ bl_int_1_24 bl_int_0_24 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c25
+ bl_int_1_25 bl_int_0_25 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c26
+ bl_int_1_26 bl_int_0_26 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c27
+ bl_int_1_27 bl_int_0_27 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c28
+ bl_int_1_28 bl_int_0_28 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c29
+ bl_int_1_29 bl_int_0_29 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c30
+ bl_int_1_30 bl_int_0_30 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c31
+ bl_int_1_31 bl_int_0_31 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c32
+ bl_int_1_32 bl_int_0_32 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c33
+ bl_int_1_33 bl_int_0_33 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c34
+ bl_int_1_34 bl_int_0_34 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c35
+ bl_int_1_35 bl_int_0_35 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c36
+ bl_int_1_36 bl_int_0_36 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c37
+ bl_int_1_37 bl_int_0_37 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c38
+ bl_int_1_38 bl_int_0_38 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c39
+ bl_int_1_39 bl_int_0_39 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c40
+ bl_int_1_40 bl_int_0_40 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c41
+ bl_int_1_41 bl_int_0_41 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c42
+ bl_int_1_42 bl_int_0_42 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c43
+ bl_int_1_43 bl_int_0_43 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c44
+ bl_int_1_44 bl_int_0_44 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c45
+ bl_int_1_45 bl_int_0_45 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c46
+ bl_int_1_46 bl_int_0_46 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c47
+ bl_int_1_47 bl_int_0_47 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c48
+ bl_int_1_48 bl_int_0_48 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c49
+ bl_int_1_49 bl_int_0_49 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c50
+ bl_int_1_50 bl_int_0_50 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c51
+ bl_int_1_51 bl_int_0_51 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c52
+ bl_int_1_52 bl_int_0_52 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c53
+ bl_int_1_53 bl_int_0_53 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c54
+ bl_int_1_54 bl_int_0_54 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c55
+ bl_int_1_55 bl_int_0_55 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c56
+ bl_int_1_56 bl_int_0_56 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c57
+ bl_int_1_57 bl_int_0_57 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c58
+ bl_int_1_58 bl_int_0_58 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c59
+ bl_int_1_59 bl_int_0_59 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c60
+ bl_int_1_60 bl_int_0_60 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c61
+ bl_int_1_61 bl_int_0_61 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c62
+ bl_int_1_62 bl_int_0_62 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c63
+ bl_int_1_63 bl_int_0_63 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c64
+ bl_int_1_64 bl_int_0_64 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c65
+ bl_int_1_65 bl_int_0_65 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c66
+ bl_int_1_66 bl_int_0_66 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c67
+ bl_int_1_67 bl_int_0_67 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c68
+ bl_int_1_68 bl_int_0_68 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c69
+ bl_int_1_69 bl_int_0_69 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c70
+ bl_int_1_70 bl_int_0_70 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c71
+ bl_int_1_71 bl_int_0_71 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c72
+ bl_int_1_72 bl_int_0_72 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c73
+ bl_int_1_73 bl_int_0_73 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c74
+ bl_int_1_74 bl_int_0_74 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c75
+ bl_int_1_75 bl_int_0_75 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c76
+ bl_int_1_76 bl_int_0_76 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c77
+ bl_int_1_77 bl_int_0_77 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c78
+ bl_int_1_78 bl_int_0_78 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c79
+ bl_int_1_79 bl_int_0_79 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c80
+ bl_int_1_80 bl_int_0_80 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c81
+ bl_int_1_81 bl_int_0_81 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c82
+ bl_int_1_82 bl_int_0_82 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c83
+ bl_int_1_83 bl_int_0_83 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c84
+ bl_int_1_84 bl_int_0_84 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c85
+ bl_int_1_85 bl_int_0_85 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c86
+ bl_int_1_86 bl_int_0_86 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c87
+ bl_int_1_87 bl_int_0_87 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c88
+ bl_int_1_88 bl_int_0_88 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c89
+ bl_int_1_89 bl_int_0_89 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c90
+ bl_int_1_90 bl_int_0_90 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c91
+ bl_int_1_91 bl_int_0_91 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c92
+ bl_int_1_92 bl_int_0_92 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c93
+ bl_int_1_93 bl_int_0_93 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c94
+ bl_int_1_94 bl_int_0_94 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c95
+ bl_int_1_95 bl_int_0_95 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c96
+ bl_int_1_96 bl_int_0_96 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c97
+ bl_int_1_97 bl_int_0_97 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c98
+ bl_int_1_98 bl_int_0_98 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c99
+ bl_int_1_99 bl_int_0_99 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c100
+ bl_int_1_100 bl_int_0_100 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c101
+ bl_int_1_101 bl_int_0_101 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c102
+ bl_int_1_102 bl_int_0_102 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c103
+ bl_int_1_103 bl_int_0_103 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c104
+ bl_int_1_104 bl_int_0_104 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c105
+ bl_int_1_105 bl_int_0_105 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c106
+ bl_int_1_106 bl_int_0_106 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c107
+ bl_int_1_107 bl_int_0_107 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c108
+ bl_int_1_108 bl_int_0_108 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c109
+ bl_int_1_109 bl_int_0_109 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c110
+ bl_int_1_110 bl_int_0_110 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c111
+ bl_int_1_111 bl_int_0_111 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c112
+ bl_int_1_112 bl_int_0_112 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c113
+ bl_int_1_113 bl_int_0_113 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c114
+ bl_int_1_114 bl_int_0_114 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c115
+ bl_int_1_115 bl_int_0_115 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c116
+ bl_int_1_116 bl_int_0_116 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c117
+ bl_int_1_117 bl_int_0_117 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c118
+ bl_int_1_118 bl_int_0_118 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c119
+ bl_int_1_119 bl_int_0_119 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c120
+ bl_int_1_120 bl_int_0_120 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c121
+ bl_int_1_121 bl_int_0_121 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c122
+ bl_int_1_122 bl_int_0_122 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c123
+ bl_int_1_123 bl_int_0_123 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c124
+ bl_int_1_124 bl_int_0_124 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c125
+ bl_int_1_125 bl_int_0_125 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c126
+ bl_int_1_126 bl_int_0_126 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c127
+ bl_int_1_127 bl_int_0_127 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c128
+ bl_int_1_128 bl_int_0_128 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c129
+ bl_int_1_129 bl_int_0_129 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c130
+ bl_int_1_130 bl_int_0_130 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c131
+ bl_int_1_131 bl_int_0_131 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c132
+ bl_int_1_132 bl_int_0_132 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c133
+ bl_int_1_133 bl_int_0_133 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c134
+ bl_int_1_134 bl_int_0_134 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c135
+ bl_int_1_135 bl_int_0_135 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c136
+ bl_int_1_136 bl_int_0_136 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c137
+ bl_int_1_137 bl_int_0_137 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c138
+ bl_int_1_138 bl_int_0_138 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c139
+ bl_int_1_139 bl_int_0_139 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c140
+ bl_int_1_140 bl_int_0_140 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c141
+ bl_int_1_141 bl_int_0_141 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c142
+ bl_int_1_142 bl_int_0_142 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c143
+ bl_int_1_143 bl_int_0_143 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c144
+ bl_int_1_144 bl_int_0_144 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c145
+ bl_int_1_145 bl_int_0_145 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c146
+ bl_int_1_146 bl_int_0_146 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c147
+ bl_int_1_147 bl_int_0_147 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c148
+ bl_int_1_148 bl_int_0_148 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c149
+ bl_int_1_149 bl_int_0_149 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c150
+ bl_int_1_150 bl_int_0_150 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c151
+ bl_int_1_151 bl_int_0_151 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c152
+ bl_int_1_152 bl_int_0_152 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c153
+ bl_int_1_153 bl_int_0_153 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c154
+ bl_int_1_154 bl_int_0_154 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c155
+ bl_int_1_155 bl_int_0_155 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c156
+ bl_int_1_156 bl_int_0_156 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c157
+ bl_int_1_157 bl_int_0_157 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c158
+ bl_int_1_158 bl_int_0_158 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c159
+ bl_int_1_159 bl_int_0_159 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c160
+ bl_int_1_160 bl_int_0_160 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c161
+ bl_int_1_161 bl_int_0_161 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c162
+ bl_int_1_162 bl_int_0_162 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c163
+ bl_int_1_163 bl_int_0_163 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c164
+ bl_int_1_164 bl_int_0_164 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c165
+ bl_int_1_165 bl_int_0_165 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c166
+ bl_int_1_166 bl_int_0_166 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c167
+ bl_int_1_167 bl_int_0_167 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c168
+ bl_int_1_168 bl_int_0_168 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c169
+ bl_int_1_169 bl_int_0_169 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c170
+ bl_int_1_170 bl_int_0_170 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c171
+ bl_int_1_171 bl_int_0_171 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c172
+ bl_int_1_172 bl_int_0_172 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c173
+ bl_int_1_173 bl_int_0_173 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c174
+ bl_int_1_174 bl_int_0_174 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c175
+ bl_int_1_175 bl_int_0_175 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c176
+ bl_int_1_176 bl_int_0_176 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c177
+ bl_int_1_177 bl_int_0_177 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c178
+ bl_int_1_178 bl_int_0_178 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c179
+ bl_int_1_179 bl_int_0_179 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c180
+ bl_int_1_180 bl_int_0_180 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c181
+ bl_int_1_181 bl_int_0_181 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c182
+ bl_int_1_182 bl_int_0_182 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r1_c183
+ bl_int_1_183 bl_int_0_183 wl_0_1 gnd
+ sram_rom_base_one_cell
Xbit_r2_c0
+ bl_int_2_0 bl_int_1_0 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c1
+ bl_int_2_1 bl_int_1_1 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c2
+ bl_int_2_2 bl_int_1_2 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c3
+ bl_int_2_3 bl_int_1_3 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c4
+ bl_int_2_4 bl_int_1_4 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c5
+ bl_int_2_5 bl_int_1_5 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c6
+ bl_int_2_6 bl_int_1_6 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c7
+ bl_int_2_7 bl_int_1_7 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c8
+ bl_int_2_8 bl_int_1_8 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c9
+ bl_int_2_9 bl_int_1_9 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c10
+ bl_int_2_10 bl_int_1_10 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c11
+ bl_int_2_11 bl_int_1_11 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c12
+ bl_int_2_12 bl_int_1_12 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c13
+ bl_int_2_13 bl_int_1_13 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c14
+ bl_int_2_14 bl_int_1_14 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c15
+ bl_int_2_15 bl_int_1_15 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c16
+ bl_int_2_16 bl_int_1_16 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c17
+ bl_int_2_17 bl_int_1_17 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c18
+ bl_int_2_18 bl_int_1_18 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c19
+ bl_int_2_19 bl_int_1_19 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c20
+ bl_int_2_20 bl_int_1_20 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c21
+ bl_int_2_21 bl_int_1_21 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c22
+ bl_int_2_22 bl_int_1_22 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c23
+ bl_int_2_23 bl_int_1_23 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c24
+ bl_int_2_24 bl_int_1_24 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c25
+ bl_int_2_25 bl_int_1_25 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c26
+ bl_int_2_26 bl_int_1_26 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c27
+ bl_int_2_27 bl_int_1_27 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c28
+ bl_int_2_28 bl_int_1_28 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c29
+ bl_int_2_29 bl_int_1_29 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c30
+ bl_int_2_30 bl_int_1_30 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c31
+ bl_int_2_31 bl_int_1_31 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c32
+ bl_int_2_32 bl_int_1_32 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c33
+ bl_int_2_33 bl_int_1_33 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c34
+ bl_int_2_34 bl_int_1_34 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c35
+ bl_int_2_35 bl_int_1_35 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c36
+ bl_int_2_36 bl_int_1_36 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c37
+ bl_int_2_37 bl_int_1_37 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c38
+ bl_int_2_38 bl_int_1_38 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c39
+ bl_int_2_39 bl_int_1_39 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c40
+ bl_int_2_40 bl_int_1_40 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c41
+ bl_int_2_41 bl_int_1_41 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c42
+ bl_int_2_42 bl_int_1_42 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c43
+ bl_int_2_43 bl_int_1_43 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c44
+ bl_int_2_44 bl_int_1_44 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c45
+ bl_int_2_45 bl_int_1_45 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c46
+ bl_int_2_46 bl_int_1_46 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c47
+ bl_int_2_47 bl_int_1_47 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c48
+ bl_int_2_48 bl_int_1_48 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c49
+ bl_int_2_49 bl_int_1_49 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c50
+ bl_int_2_50 bl_int_1_50 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c51
+ bl_int_2_51 bl_int_1_51 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c52
+ bl_int_2_52 bl_int_1_52 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c53
+ bl_int_2_53 bl_int_1_53 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c54
+ bl_int_2_54 bl_int_1_54 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c55
+ bl_int_2_55 bl_int_1_55 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c56
+ bl_int_2_56 bl_int_1_56 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c57
+ bl_int_2_57 bl_int_1_57 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c58
+ bl_int_2_58 bl_int_1_58 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c59
+ bl_int_2_59 bl_int_1_59 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c60
+ bl_int_2_60 bl_int_1_60 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c61
+ bl_int_2_61 bl_int_1_61 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c62
+ bl_int_2_62 bl_int_1_62 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c63
+ bl_int_2_63 bl_int_1_63 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c64
+ bl_int_2_64 bl_int_1_64 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c65
+ bl_int_2_65 bl_int_1_65 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c66
+ bl_int_2_66 bl_int_1_66 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c67
+ bl_int_2_67 bl_int_1_67 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c68
+ bl_int_2_68 bl_int_1_68 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c69
+ bl_int_2_69 bl_int_1_69 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c70
+ bl_int_2_70 bl_int_1_70 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c71
+ bl_int_2_71 bl_int_1_71 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c72
+ bl_int_2_72 bl_int_1_72 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c73
+ bl_int_2_73 bl_int_1_73 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c74
+ bl_int_2_74 bl_int_1_74 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c75
+ bl_int_2_75 bl_int_1_75 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c76
+ bl_int_2_76 bl_int_1_76 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c77
+ bl_int_2_77 bl_int_1_77 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c78
+ bl_int_2_78 bl_int_1_78 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c79
+ bl_int_2_79 bl_int_1_79 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c80
+ bl_int_2_80 bl_int_1_80 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c81
+ bl_int_2_81 bl_int_1_81 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c82
+ bl_int_2_82 bl_int_1_82 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c83
+ bl_int_2_83 bl_int_1_83 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c84
+ bl_int_2_84 bl_int_1_84 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c85
+ bl_int_2_85 bl_int_1_85 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c86
+ bl_int_2_86 bl_int_1_86 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c87
+ bl_int_2_87 bl_int_1_87 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c88
+ bl_int_2_88 bl_int_1_88 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c89
+ bl_int_2_89 bl_int_1_89 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c90
+ bl_int_2_90 bl_int_1_90 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c91
+ bl_int_2_91 bl_int_1_91 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c92
+ bl_int_2_92 bl_int_1_92 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c93
+ bl_int_2_93 bl_int_1_93 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c94
+ bl_int_2_94 bl_int_1_94 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c95
+ bl_int_2_95 bl_int_1_95 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c96
+ bl_int_2_96 bl_int_1_96 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c97
+ bl_int_2_97 bl_int_1_97 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c98
+ bl_int_2_98 bl_int_1_98 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c99
+ bl_int_2_99 bl_int_1_99 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c100
+ bl_int_2_100 bl_int_1_100 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c101
+ bl_int_2_101 bl_int_1_101 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c102
+ bl_int_2_102 bl_int_1_102 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c103
+ bl_int_2_103 bl_int_1_103 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c104
+ bl_int_2_104 bl_int_1_104 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c105
+ bl_int_2_105 bl_int_1_105 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c106
+ bl_int_2_106 bl_int_1_106 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c107
+ bl_int_2_107 bl_int_1_107 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c108
+ bl_int_2_108 bl_int_1_108 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c109
+ bl_int_2_109 bl_int_1_109 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c110
+ bl_int_2_110 bl_int_1_110 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c111
+ bl_int_2_111 bl_int_1_111 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c112
+ bl_int_2_112 bl_int_1_112 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c113
+ bl_int_2_113 bl_int_1_113 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c114
+ bl_int_2_114 bl_int_1_114 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c115
+ bl_int_2_115 bl_int_1_115 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c116
+ bl_int_2_116 bl_int_1_116 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c117
+ bl_int_2_117 bl_int_1_117 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c118
+ bl_int_2_118 bl_int_1_118 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c119
+ bl_int_2_119 bl_int_1_119 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c120
+ bl_int_2_120 bl_int_1_120 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c121
+ bl_int_2_121 bl_int_1_121 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c122
+ bl_int_2_122 bl_int_1_122 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c123
+ bl_int_2_123 bl_int_1_123 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c124
+ bl_int_2_124 bl_int_1_124 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c125
+ bl_int_2_125 bl_int_1_125 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c126
+ bl_int_2_126 bl_int_1_126 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c127
+ bl_int_2_127 bl_int_1_127 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c128
+ bl_int_2_128 bl_int_1_128 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c129
+ bl_int_2_129 bl_int_1_129 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c130
+ bl_int_2_130 bl_int_1_130 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c131
+ bl_int_2_131 bl_int_1_131 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c132
+ bl_int_2_132 bl_int_1_132 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c133
+ bl_int_2_133 bl_int_1_133 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c134
+ bl_int_2_134 bl_int_1_134 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c135
+ bl_int_2_135 bl_int_1_135 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c136
+ bl_int_2_136 bl_int_1_136 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c137
+ bl_int_2_137 bl_int_1_137 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c138
+ bl_int_2_138 bl_int_1_138 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c139
+ bl_int_2_139 bl_int_1_139 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c140
+ bl_int_2_140 bl_int_1_140 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c141
+ bl_int_2_141 bl_int_1_141 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c142
+ bl_int_2_142 bl_int_1_142 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c143
+ bl_int_2_143 bl_int_1_143 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c144
+ bl_int_2_144 bl_int_1_144 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c145
+ bl_int_2_145 bl_int_1_145 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c146
+ bl_int_2_146 bl_int_1_146 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c147
+ bl_int_2_147 bl_int_1_147 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c148
+ bl_int_2_148 bl_int_1_148 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c149
+ bl_int_2_149 bl_int_1_149 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c150
+ bl_int_2_150 bl_int_1_150 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c151
+ bl_int_2_151 bl_int_1_151 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c152
+ bl_int_2_152 bl_int_1_152 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c153
+ bl_int_2_153 bl_int_1_153 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c154
+ bl_int_2_154 bl_int_1_154 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c155
+ bl_int_2_155 bl_int_1_155 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c156
+ bl_int_2_156 bl_int_1_156 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c157
+ bl_int_2_157 bl_int_1_157 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c158
+ bl_int_2_158 bl_int_1_158 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c159
+ bl_int_2_159 bl_int_1_159 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c160
+ bl_int_2_160 bl_int_1_160 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c161
+ bl_int_2_161 bl_int_1_161 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c162
+ bl_int_2_162 bl_int_1_162 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c163
+ bl_int_2_163 bl_int_1_163 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c164
+ bl_int_2_164 bl_int_1_164 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c165
+ bl_int_2_165 bl_int_1_165 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c166
+ bl_int_2_166 bl_int_1_166 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c167
+ bl_int_2_167 bl_int_1_167 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c168
+ bl_int_2_168 bl_int_1_168 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c169
+ bl_int_2_169 bl_int_1_169 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c170
+ bl_int_2_170 bl_int_1_170 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c171
+ bl_int_2_171 bl_int_1_171 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c172
+ bl_int_2_172 bl_int_1_172 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c173
+ bl_int_2_173 bl_int_1_173 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c174
+ bl_int_2_174 bl_int_1_174 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c175
+ bl_int_2_175 bl_int_1_175 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c176
+ bl_int_2_176 bl_int_1_176 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c177
+ bl_int_2_177 bl_int_1_177 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c178
+ bl_int_2_178 bl_int_1_178 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c179
+ bl_int_2_179 bl_int_1_179 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c180
+ bl_int_2_180 bl_int_1_180 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c181
+ bl_int_2_181 bl_int_1_181 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c182
+ bl_int_2_182 bl_int_1_182 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r2_c183
+ bl_int_2_183 bl_int_1_183 wl_0_2 gnd
+ sram_rom_base_one_cell
Xbit_r3_c0
+ bl_int_3_0 bl_int_2_0 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c1
+ bl_int_3_1 bl_int_2_1 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c2
+ bl_int_3_2 bl_int_2_2 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c3
+ bl_int_3_3 bl_int_2_3 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c4
+ bl_int_3_4 bl_int_2_4 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c5
+ bl_int_3_5 bl_int_2_5 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c6
+ bl_int_3_6 bl_int_2_6 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c7
+ bl_int_3_7 bl_int_2_7 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c8
+ bl_int_3_8 bl_int_2_8 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c9
+ bl_int_3_9 bl_int_2_9 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c10
+ bl_int_3_10 bl_int_2_10 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c11
+ bl_int_3_11 bl_int_2_11 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c12
+ bl_int_3_12 bl_int_2_12 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c13
+ bl_int_3_13 bl_int_2_13 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c14
+ bl_int_3_14 bl_int_2_14 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c15
+ bl_int_3_15 bl_int_2_15 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c16
+ bl_int_3_16 bl_int_2_16 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c17
+ bl_int_3_17 bl_int_2_17 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c18
+ bl_int_3_18 bl_int_2_18 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c19
+ bl_int_3_19 bl_int_2_19 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c20
+ bl_int_3_20 bl_int_2_20 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c21
+ bl_int_3_21 bl_int_2_21 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c22
+ bl_int_3_22 bl_int_2_22 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c23
+ bl_int_3_23 bl_int_2_23 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c24
+ bl_int_3_24 bl_int_2_24 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c25
+ bl_int_3_25 bl_int_2_25 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c26
+ bl_int_3_26 bl_int_2_26 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c27
+ bl_int_3_27 bl_int_2_27 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c28
+ bl_int_3_28 bl_int_2_28 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c29
+ bl_int_3_29 bl_int_2_29 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c30
+ bl_int_3_30 bl_int_2_30 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c31
+ bl_int_3_31 bl_int_2_31 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c32
+ bl_int_3_32 bl_int_2_32 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c33
+ bl_int_3_33 bl_int_2_33 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c34
+ bl_int_3_34 bl_int_2_34 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c35
+ bl_int_3_35 bl_int_2_35 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c36
+ bl_int_3_36 bl_int_2_36 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c37
+ bl_int_3_37 bl_int_2_37 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c38
+ bl_int_3_38 bl_int_2_38 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c39
+ bl_int_3_39 bl_int_2_39 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c40
+ bl_int_3_40 bl_int_2_40 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c41
+ bl_int_3_41 bl_int_2_41 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c42
+ bl_int_3_42 bl_int_2_42 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c43
+ bl_int_3_43 bl_int_2_43 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c44
+ bl_int_3_44 bl_int_2_44 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c45
+ bl_int_3_45 bl_int_2_45 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c46
+ bl_int_3_46 bl_int_2_46 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c47
+ bl_int_3_47 bl_int_2_47 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c48
+ bl_int_3_48 bl_int_2_48 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c49
+ bl_int_3_49 bl_int_2_49 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c50
+ bl_int_3_50 bl_int_2_50 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c51
+ bl_int_3_51 bl_int_2_51 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c52
+ bl_int_3_52 bl_int_2_52 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c53
+ bl_int_3_53 bl_int_2_53 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c54
+ bl_int_3_54 bl_int_2_54 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c55
+ bl_int_3_55 bl_int_2_55 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c56
+ bl_int_3_56 bl_int_2_56 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c57
+ bl_int_3_57 bl_int_2_57 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c58
+ bl_int_3_58 bl_int_2_58 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c59
+ bl_int_3_59 bl_int_2_59 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c60
+ bl_int_3_60 bl_int_2_60 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c61
+ bl_int_3_61 bl_int_2_61 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c62
+ bl_int_3_62 bl_int_2_62 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c63
+ bl_int_3_63 bl_int_2_63 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c64
+ bl_int_3_64 bl_int_2_64 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c65
+ bl_int_3_65 bl_int_2_65 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c66
+ bl_int_3_66 bl_int_2_66 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c67
+ bl_int_3_67 bl_int_2_67 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c68
+ bl_int_3_68 bl_int_2_68 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c69
+ bl_int_3_69 bl_int_2_69 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c70
+ bl_int_3_70 bl_int_2_70 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c71
+ bl_int_3_71 bl_int_2_71 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c72
+ bl_int_3_72 bl_int_2_72 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c73
+ bl_int_3_73 bl_int_2_73 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c74
+ bl_int_3_74 bl_int_2_74 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c75
+ bl_int_3_75 bl_int_2_75 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c76
+ bl_int_3_76 bl_int_2_76 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c77
+ bl_int_3_77 bl_int_2_77 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c78
+ bl_int_3_78 bl_int_2_78 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c79
+ bl_int_3_79 bl_int_2_79 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c80
+ bl_int_3_80 bl_int_2_80 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c81
+ bl_int_3_81 bl_int_2_81 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c82
+ bl_int_3_82 bl_int_2_82 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c83
+ bl_int_3_83 bl_int_2_83 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c84
+ bl_int_3_84 bl_int_2_84 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c85
+ bl_int_3_85 bl_int_2_85 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c86
+ bl_int_3_86 bl_int_2_86 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c87
+ bl_int_3_87 bl_int_2_87 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c88
+ bl_int_3_88 bl_int_2_88 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c89
+ bl_int_3_89 bl_int_2_89 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c90
+ bl_int_3_90 bl_int_2_90 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c91
+ bl_int_3_91 bl_int_2_91 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c92
+ bl_int_3_92 bl_int_2_92 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c93
+ bl_int_3_93 bl_int_2_93 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c94
+ bl_int_3_94 bl_int_2_94 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c95
+ bl_int_3_95 bl_int_2_95 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c96
+ bl_int_3_96 bl_int_2_96 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c97
+ bl_int_3_97 bl_int_2_97 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c98
+ bl_int_3_98 bl_int_2_98 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c99
+ bl_int_3_99 bl_int_2_99 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c100
+ bl_int_3_100 bl_int_2_100 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c101
+ bl_int_3_101 bl_int_2_101 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c102
+ bl_int_3_102 bl_int_2_102 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c103
+ bl_int_3_103 bl_int_2_103 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c104
+ bl_int_3_104 bl_int_2_104 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c105
+ bl_int_3_105 bl_int_2_105 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c106
+ bl_int_3_106 bl_int_2_106 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c107
+ bl_int_3_107 bl_int_2_107 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c108
+ bl_int_3_108 bl_int_2_108 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c109
+ bl_int_3_109 bl_int_2_109 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c110
+ bl_int_3_110 bl_int_2_110 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c111
+ bl_int_3_111 bl_int_2_111 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c112
+ bl_int_3_112 bl_int_2_112 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c113
+ bl_int_3_113 bl_int_2_113 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c114
+ bl_int_3_114 bl_int_2_114 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c115
+ bl_int_3_115 bl_int_2_115 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c116
+ bl_int_3_116 bl_int_2_116 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c117
+ bl_int_3_117 bl_int_2_117 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c118
+ bl_int_3_118 bl_int_2_118 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c119
+ bl_int_3_119 bl_int_2_119 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c120
+ bl_int_3_120 bl_int_2_120 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c121
+ bl_int_3_121 bl_int_2_121 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c122
+ bl_int_3_122 bl_int_2_122 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c123
+ bl_int_3_123 bl_int_2_123 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c124
+ bl_int_3_124 bl_int_2_124 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c125
+ bl_int_3_125 bl_int_2_125 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c126
+ bl_int_3_126 bl_int_2_126 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c127
+ bl_int_3_127 bl_int_2_127 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c128
+ bl_int_3_128 bl_int_2_128 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c129
+ bl_int_3_129 bl_int_2_129 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c130
+ bl_int_3_130 bl_int_2_130 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c131
+ bl_int_3_131 bl_int_2_131 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c132
+ bl_int_3_132 bl_int_2_132 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c133
+ bl_int_3_133 bl_int_2_133 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c134
+ bl_int_3_134 bl_int_2_134 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c135
+ bl_int_3_135 bl_int_2_135 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c136
+ bl_int_3_136 bl_int_2_136 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c137
+ bl_int_3_137 bl_int_2_137 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c138
+ bl_int_3_138 bl_int_2_138 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c139
+ bl_int_3_139 bl_int_2_139 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c140
+ bl_int_3_140 bl_int_2_140 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c141
+ bl_int_3_141 bl_int_2_141 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c142
+ bl_int_3_142 bl_int_2_142 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c143
+ bl_int_3_143 bl_int_2_143 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c144
+ bl_int_3_144 bl_int_2_144 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c145
+ bl_int_3_145 bl_int_2_145 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c146
+ bl_int_3_146 bl_int_2_146 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c147
+ bl_int_3_147 bl_int_2_147 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c148
+ bl_int_3_148 bl_int_2_148 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c149
+ bl_int_3_149 bl_int_2_149 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c150
+ bl_int_3_150 bl_int_2_150 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c151
+ bl_int_3_151 bl_int_2_151 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c152
+ bl_int_3_152 bl_int_2_152 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c153
+ bl_int_3_153 bl_int_2_153 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c154
+ bl_int_3_154 bl_int_2_154 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c155
+ bl_int_3_155 bl_int_2_155 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c156
+ bl_int_3_156 bl_int_2_156 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c157
+ bl_int_3_157 bl_int_2_157 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c158
+ bl_int_3_158 bl_int_2_158 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c159
+ bl_int_3_159 bl_int_2_159 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c160
+ bl_int_3_160 bl_int_2_160 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c161
+ bl_int_3_161 bl_int_2_161 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c162
+ bl_int_3_162 bl_int_2_162 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c163
+ bl_int_3_163 bl_int_2_163 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c164
+ bl_int_3_164 bl_int_2_164 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c165
+ bl_int_3_165 bl_int_2_165 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c166
+ bl_int_3_166 bl_int_2_166 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c167
+ bl_int_3_167 bl_int_2_167 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c168
+ bl_int_3_168 bl_int_2_168 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c169
+ bl_int_3_169 bl_int_2_169 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c170
+ bl_int_3_170 bl_int_2_170 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c171
+ bl_int_3_171 bl_int_2_171 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c172
+ bl_int_3_172 bl_int_2_172 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c173
+ bl_int_3_173 bl_int_2_173 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c174
+ bl_int_3_174 bl_int_2_174 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c175
+ bl_int_3_175 bl_int_2_175 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c176
+ bl_int_3_176 bl_int_2_176 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c177
+ bl_int_3_177 bl_int_2_177 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c178
+ bl_int_3_178 bl_int_2_178 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c179
+ bl_int_3_179 bl_int_2_179 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c180
+ bl_int_3_180 bl_int_2_180 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c181
+ bl_int_3_181 bl_int_2_181 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c182
+ bl_int_3_182 bl_int_2_182 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r3_c183
+ bl_int_3_183 bl_int_2_183 wl_0_3 gnd
+ sram_rom_base_one_cell
Xbit_r4_c0
+ bl_int_4_0 bl_int_3_0 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c1
+ bl_int_4_1 bl_int_3_1 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c2
+ bl_int_4_2 bl_int_3_2 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c3
+ bl_int_4_3 bl_int_3_3 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c4
+ bl_int_4_4 bl_int_3_4 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c5
+ bl_int_4_5 bl_int_3_5 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c6
+ bl_int_4_6 bl_int_3_6 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c7
+ bl_int_4_7 bl_int_3_7 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c8
+ bl_int_4_8 bl_int_3_8 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c9
+ bl_int_4_9 bl_int_3_9 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c10
+ bl_int_4_10 bl_int_3_10 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c11
+ bl_int_4_11 bl_int_3_11 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c12
+ bl_int_4_12 bl_int_3_12 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c13
+ bl_int_4_13 bl_int_3_13 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c14
+ bl_int_4_14 bl_int_3_14 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c15
+ bl_int_4_15 bl_int_3_15 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c16
+ bl_int_4_16 bl_int_3_16 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c17
+ bl_int_4_17 bl_int_3_17 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c18
+ bl_int_4_18 bl_int_3_18 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c19
+ bl_int_4_19 bl_int_3_19 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c20
+ bl_int_4_20 bl_int_3_20 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c21
+ bl_int_4_21 bl_int_3_21 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c22
+ bl_int_4_22 bl_int_3_22 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c23
+ bl_int_4_23 bl_int_3_23 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c24
+ bl_int_4_24 bl_int_3_24 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c25
+ bl_int_4_25 bl_int_3_25 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c26
+ bl_int_4_26 bl_int_3_26 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c27
+ bl_int_4_27 bl_int_3_27 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c28
+ bl_int_4_28 bl_int_3_28 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c29
+ bl_int_4_29 bl_int_3_29 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c30
+ bl_int_4_30 bl_int_3_30 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c31
+ bl_int_4_31 bl_int_3_31 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c32
+ bl_int_4_32 bl_int_3_32 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c33
+ bl_int_4_33 bl_int_3_33 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c34
+ bl_int_4_34 bl_int_3_34 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c35
+ bl_int_4_35 bl_int_3_35 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c36
+ bl_int_4_36 bl_int_3_36 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c37
+ bl_int_4_37 bl_int_3_37 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c38
+ bl_int_4_38 bl_int_3_38 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c39
+ bl_int_4_39 bl_int_3_39 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c40
+ bl_int_4_40 bl_int_3_40 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c41
+ bl_int_4_41 bl_int_3_41 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c42
+ bl_int_4_42 bl_int_3_42 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c43
+ bl_int_4_43 bl_int_3_43 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c44
+ bl_int_4_44 bl_int_3_44 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c45
+ bl_int_4_45 bl_int_3_45 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c46
+ bl_int_4_46 bl_int_3_46 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c47
+ bl_int_4_47 bl_int_3_47 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c48
+ bl_int_4_48 bl_int_3_48 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c49
+ bl_int_4_49 bl_int_3_49 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c50
+ bl_int_4_50 bl_int_3_50 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c51
+ bl_int_4_51 bl_int_3_51 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c52
+ bl_int_4_52 bl_int_3_52 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c53
+ bl_int_4_53 bl_int_3_53 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c54
+ bl_int_4_54 bl_int_3_54 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c55
+ bl_int_4_55 bl_int_3_55 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c56
+ bl_int_4_56 bl_int_3_56 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c57
+ bl_int_4_57 bl_int_3_57 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c58
+ bl_int_4_58 bl_int_3_58 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c59
+ bl_int_4_59 bl_int_3_59 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c60
+ bl_int_4_60 bl_int_3_60 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c61
+ bl_int_4_61 bl_int_3_61 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c62
+ bl_int_4_62 bl_int_3_62 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c63
+ bl_int_4_63 bl_int_3_63 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c64
+ bl_int_4_64 bl_int_3_64 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c65
+ bl_int_4_65 bl_int_3_65 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c66
+ bl_int_4_66 bl_int_3_66 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c67
+ bl_int_4_67 bl_int_3_67 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c68
+ bl_int_4_68 bl_int_3_68 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c69
+ bl_int_4_69 bl_int_3_69 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c70
+ bl_int_4_70 bl_int_3_70 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c71
+ bl_int_4_71 bl_int_3_71 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c72
+ bl_int_4_72 bl_int_3_72 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c73
+ bl_int_4_73 bl_int_3_73 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c74
+ bl_int_4_74 bl_int_3_74 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c75
+ bl_int_4_75 bl_int_3_75 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c76
+ bl_int_4_76 bl_int_3_76 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c77
+ bl_int_4_77 bl_int_3_77 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c78
+ bl_int_4_78 bl_int_3_78 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c79
+ bl_int_4_79 bl_int_3_79 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c80
+ bl_int_4_80 bl_int_3_80 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c81
+ bl_int_4_81 bl_int_3_81 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c82
+ bl_int_4_82 bl_int_3_82 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c83
+ bl_int_4_83 bl_int_3_83 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c84
+ bl_int_4_84 bl_int_3_84 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c85
+ bl_int_4_85 bl_int_3_85 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c86
+ bl_int_4_86 bl_int_3_86 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c87
+ bl_int_4_87 bl_int_3_87 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c88
+ bl_int_4_88 bl_int_3_88 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c89
+ bl_int_4_89 bl_int_3_89 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c90
+ bl_int_4_90 bl_int_3_90 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c91
+ bl_int_4_91 bl_int_3_91 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c92
+ bl_int_4_92 bl_int_3_92 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c93
+ bl_int_4_93 bl_int_3_93 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c94
+ bl_int_4_94 bl_int_3_94 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c95
+ bl_int_4_95 bl_int_3_95 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c96
+ bl_int_4_96 bl_int_3_96 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c97
+ bl_int_4_97 bl_int_3_97 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c98
+ bl_int_4_98 bl_int_3_98 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c99
+ bl_int_4_99 bl_int_3_99 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c100
+ bl_int_4_100 bl_int_3_100 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c101
+ bl_int_4_101 bl_int_3_101 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c102
+ bl_int_4_102 bl_int_3_102 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c103
+ bl_int_4_103 bl_int_3_103 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c104
+ bl_int_4_104 bl_int_3_104 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c105
+ bl_int_4_105 bl_int_3_105 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c106
+ bl_int_4_106 bl_int_3_106 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c107
+ bl_int_4_107 bl_int_3_107 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c108
+ bl_int_4_108 bl_int_3_108 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c109
+ bl_int_4_109 bl_int_3_109 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c110
+ bl_int_4_110 bl_int_3_110 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c111
+ bl_int_4_111 bl_int_3_111 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c112
+ bl_int_4_112 bl_int_3_112 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c113
+ bl_int_4_113 bl_int_3_113 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c114
+ bl_int_4_114 bl_int_3_114 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c115
+ bl_int_4_115 bl_int_3_115 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c116
+ bl_int_4_116 bl_int_3_116 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c117
+ bl_int_4_117 bl_int_3_117 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c118
+ bl_int_4_118 bl_int_3_118 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c119
+ bl_int_4_119 bl_int_3_119 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c120
+ bl_int_4_120 bl_int_3_120 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c121
+ bl_int_4_121 bl_int_3_121 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c122
+ bl_int_4_122 bl_int_3_122 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c123
+ bl_int_4_123 bl_int_3_123 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c124
+ bl_int_4_124 bl_int_3_124 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c125
+ bl_int_4_125 bl_int_3_125 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c126
+ bl_int_4_126 bl_int_3_126 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c127
+ bl_int_4_127 bl_int_3_127 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c128
+ bl_int_4_128 bl_int_3_128 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c129
+ bl_int_4_129 bl_int_3_129 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c130
+ bl_int_4_130 bl_int_3_130 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c131
+ bl_int_4_131 bl_int_3_131 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c132
+ bl_int_4_132 bl_int_3_132 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c133
+ bl_int_4_133 bl_int_3_133 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c134
+ bl_int_4_134 bl_int_3_134 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c135
+ bl_int_4_135 bl_int_3_135 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c136
+ bl_int_4_136 bl_int_3_136 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c137
+ bl_int_4_137 bl_int_3_137 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c138
+ bl_int_4_138 bl_int_3_138 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c139
+ bl_int_4_139 bl_int_3_139 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c140
+ bl_int_4_140 bl_int_3_140 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c141
+ bl_int_4_141 bl_int_3_141 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c142
+ bl_int_4_142 bl_int_3_142 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c143
+ bl_int_4_143 bl_int_3_143 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c144
+ bl_int_4_144 bl_int_3_144 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c145
+ bl_int_4_145 bl_int_3_145 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c146
+ bl_int_4_146 bl_int_3_146 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c147
+ bl_int_4_147 bl_int_3_147 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c148
+ bl_int_4_148 bl_int_3_148 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c149
+ bl_int_4_149 bl_int_3_149 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c150
+ bl_int_4_150 bl_int_3_150 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c151
+ bl_int_4_151 bl_int_3_151 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c152
+ bl_int_4_152 bl_int_3_152 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c153
+ bl_int_4_153 bl_int_3_153 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c154
+ bl_int_4_154 bl_int_3_154 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c155
+ bl_int_4_155 bl_int_3_155 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c156
+ bl_int_4_156 bl_int_3_156 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c157
+ bl_int_4_157 bl_int_3_157 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c158
+ bl_int_4_158 bl_int_3_158 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c159
+ bl_int_4_159 bl_int_3_159 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c160
+ bl_int_4_160 bl_int_3_160 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c161
+ bl_int_4_161 bl_int_3_161 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c162
+ bl_int_4_162 bl_int_3_162 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c163
+ bl_int_4_163 bl_int_3_163 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c164
+ bl_int_4_164 bl_int_3_164 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c165
+ bl_int_4_165 bl_int_3_165 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c166
+ bl_int_4_166 bl_int_3_166 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c167
+ bl_int_4_167 bl_int_3_167 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c168
+ bl_int_4_168 bl_int_3_168 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c169
+ bl_int_4_169 bl_int_3_169 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c170
+ bl_int_4_170 bl_int_3_170 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c171
+ bl_int_4_171 bl_int_3_171 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c172
+ bl_int_4_172 bl_int_3_172 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c173
+ bl_int_4_173 bl_int_3_173 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c174
+ bl_int_4_174 bl_int_3_174 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c175
+ bl_int_4_175 bl_int_3_175 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c176
+ bl_int_4_176 bl_int_3_176 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c177
+ bl_int_4_177 bl_int_3_177 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c178
+ bl_int_4_178 bl_int_3_178 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c179
+ bl_int_4_179 bl_int_3_179 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c180
+ bl_int_4_180 bl_int_3_180 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c181
+ bl_int_4_181 bl_int_3_181 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c182
+ bl_int_4_182 bl_int_3_182 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r4_c183
+ bl_int_4_183 bl_int_3_183 wl_0_4 gnd
+ sram_rom_base_one_cell
Xbit_r5_c0
+ bl_int_5_0 bl_int_4_0 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c1
+ bl_int_5_1 bl_int_4_1 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c2
+ bl_int_5_2 bl_int_4_2 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c3
+ bl_int_5_3 bl_int_4_3 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c4
+ bl_int_5_4 bl_int_4_4 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c5
+ bl_int_5_5 bl_int_4_5 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c6
+ bl_int_5_6 bl_int_4_6 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c7
+ bl_int_5_7 bl_int_4_7 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c8
+ bl_int_5_8 bl_int_4_8 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c9
+ bl_int_5_9 bl_int_4_9 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c10
+ bl_int_5_10 bl_int_4_10 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c11
+ bl_int_5_11 bl_int_4_11 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c12
+ bl_int_5_12 bl_int_4_12 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c13
+ bl_int_5_13 bl_int_4_13 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c14
+ bl_int_5_14 bl_int_4_14 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c15
+ bl_int_5_15 bl_int_4_15 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c16
+ bl_int_5_16 bl_int_4_16 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c17
+ bl_int_5_17 bl_int_4_17 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c18
+ bl_int_5_18 bl_int_4_18 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c19
+ bl_int_5_19 bl_int_4_19 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c20
+ bl_int_5_20 bl_int_4_20 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c21
+ bl_int_5_21 bl_int_4_21 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c22
+ bl_int_5_22 bl_int_4_22 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c23
+ bl_int_5_23 bl_int_4_23 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c24
+ bl_int_5_24 bl_int_4_24 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c25
+ bl_int_5_25 bl_int_4_25 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c26
+ bl_int_5_26 bl_int_4_26 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c27
+ bl_int_5_27 bl_int_4_27 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c28
+ bl_int_5_28 bl_int_4_28 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c29
+ bl_int_5_29 bl_int_4_29 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c30
+ bl_int_5_30 bl_int_4_30 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c31
+ bl_int_5_31 bl_int_4_31 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c32
+ bl_int_5_32 bl_int_4_32 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c33
+ bl_int_5_33 bl_int_4_33 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c34
+ bl_int_5_34 bl_int_4_34 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c35
+ bl_int_5_35 bl_int_4_35 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c36
+ bl_int_5_36 bl_int_4_36 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c37
+ bl_int_5_37 bl_int_4_37 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c38
+ bl_int_5_38 bl_int_4_38 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c39
+ bl_int_5_39 bl_int_4_39 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c40
+ bl_int_5_40 bl_int_4_40 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c41
+ bl_int_5_41 bl_int_4_41 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c42
+ bl_int_5_42 bl_int_4_42 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c43
+ bl_int_5_43 bl_int_4_43 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c44
+ bl_int_5_44 bl_int_4_44 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c45
+ bl_int_5_45 bl_int_4_45 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c46
+ bl_int_5_46 bl_int_4_46 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c47
+ bl_int_5_47 bl_int_4_47 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c48
+ bl_int_5_48 bl_int_4_48 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c49
+ bl_int_5_49 bl_int_4_49 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c50
+ bl_int_5_50 bl_int_4_50 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c51
+ bl_int_5_51 bl_int_4_51 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c52
+ bl_int_5_52 bl_int_4_52 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c53
+ bl_int_5_53 bl_int_4_53 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c54
+ bl_int_5_54 bl_int_4_54 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c55
+ bl_int_5_55 bl_int_4_55 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c56
+ bl_int_5_56 bl_int_4_56 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c57
+ bl_int_5_57 bl_int_4_57 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c58
+ bl_int_5_58 bl_int_4_58 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c59
+ bl_int_5_59 bl_int_4_59 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c60
+ bl_int_5_60 bl_int_4_60 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c61
+ bl_int_5_61 bl_int_4_61 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c62
+ bl_int_5_62 bl_int_4_62 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c63
+ bl_int_5_63 bl_int_4_63 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c64
+ bl_int_5_64 bl_int_4_64 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c65
+ bl_int_5_65 bl_int_4_65 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c66
+ bl_int_5_66 bl_int_4_66 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c67
+ bl_int_5_67 bl_int_4_67 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c68
+ bl_int_5_68 bl_int_4_68 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c69
+ bl_int_5_69 bl_int_4_69 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c70
+ bl_int_5_70 bl_int_4_70 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c71
+ bl_int_5_71 bl_int_4_71 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c72
+ bl_int_5_72 bl_int_4_72 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c73
+ bl_int_5_73 bl_int_4_73 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c74
+ bl_int_5_74 bl_int_4_74 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c75
+ bl_int_5_75 bl_int_4_75 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c76
+ bl_int_5_76 bl_int_4_76 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c77
+ bl_int_5_77 bl_int_4_77 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c78
+ bl_int_5_78 bl_int_4_78 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c79
+ bl_int_5_79 bl_int_4_79 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c80
+ bl_int_5_80 bl_int_4_80 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c81
+ bl_int_5_81 bl_int_4_81 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c82
+ bl_int_5_82 bl_int_4_82 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c83
+ bl_int_5_83 bl_int_4_83 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c84
+ bl_int_5_84 bl_int_4_84 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c85
+ bl_int_5_85 bl_int_4_85 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c86
+ bl_int_5_86 bl_int_4_86 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c87
+ bl_int_5_87 bl_int_4_87 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c88
+ bl_int_5_88 bl_int_4_88 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c89
+ bl_int_5_89 bl_int_4_89 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c90
+ bl_int_5_90 bl_int_4_90 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c91
+ bl_int_5_91 bl_int_4_91 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c92
+ bl_int_5_92 bl_int_4_92 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c93
+ bl_int_5_93 bl_int_4_93 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c94
+ bl_int_5_94 bl_int_4_94 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c95
+ bl_int_5_95 bl_int_4_95 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c96
+ bl_int_5_96 bl_int_4_96 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c97
+ bl_int_5_97 bl_int_4_97 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c98
+ bl_int_5_98 bl_int_4_98 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c99
+ bl_int_5_99 bl_int_4_99 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c100
+ bl_int_5_100 bl_int_4_100 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c101
+ bl_int_5_101 bl_int_4_101 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c102
+ bl_int_5_102 bl_int_4_102 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c103
+ bl_int_5_103 bl_int_4_103 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c104
+ bl_int_5_104 bl_int_4_104 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c105
+ bl_int_5_105 bl_int_4_105 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c106
+ bl_int_5_106 bl_int_4_106 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c107
+ bl_int_5_107 bl_int_4_107 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c108
+ bl_int_5_108 bl_int_4_108 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c109
+ bl_int_5_109 bl_int_4_109 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c110
+ bl_int_5_110 bl_int_4_110 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c111
+ bl_int_5_111 bl_int_4_111 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c112
+ bl_int_5_112 bl_int_4_112 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c113
+ bl_int_5_113 bl_int_4_113 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c114
+ bl_int_5_114 bl_int_4_114 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c115
+ bl_int_5_115 bl_int_4_115 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c116
+ bl_int_5_116 bl_int_4_116 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c117
+ bl_int_5_117 bl_int_4_117 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c118
+ bl_int_5_118 bl_int_4_118 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c119
+ bl_int_5_119 bl_int_4_119 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c120
+ bl_int_5_120 bl_int_4_120 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c121
+ bl_int_5_121 bl_int_4_121 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c122
+ bl_int_5_122 bl_int_4_122 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c123
+ bl_int_5_123 bl_int_4_123 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c124
+ bl_int_5_124 bl_int_4_124 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c125
+ bl_int_5_125 bl_int_4_125 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c126
+ bl_int_5_126 bl_int_4_126 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c127
+ bl_int_5_127 bl_int_4_127 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c128
+ bl_int_5_128 bl_int_4_128 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c129
+ bl_int_5_129 bl_int_4_129 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c130
+ bl_int_5_130 bl_int_4_130 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c131
+ bl_int_5_131 bl_int_4_131 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c132
+ bl_int_5_132 bl_int_4_132 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c133
+ bl_int_5_133 bl_int_4_133 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c134
+ bl_int_5_134 bl_int_4_134 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c135
+ bl_int_5_135 bl_int_4_135 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c136
+ bl_int_5_136 bl_int_4_136 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c137
+ bl_int_5_137 bl_int_4_137 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c138
+ bl_int_5_138 bl_int_4_138 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c139
+ bl_int_5_139 bl_int_4_139 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c140
+ bl_int_5_140 bl_int_4_140 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c141
+ bl_int_5_141 bl_int_4_141 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c142
+ bl_int_5_142 bl_int_4_142 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c143
+ bl_int_5_143 bl_int_4_143 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c144
+ bl_int_5_144 bl_int_4_144 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c145
+ bl_int_5_145 bl_int_4_145 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c146
+ bl_int_5_146 bl_int_4_146 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c147
+ bl_int_5_147 bl_int_4_147 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c148
+ bl_int_5_148 bl_int_4_148 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c149
+ bl_int_5_149 bl_int_4_149 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c150
+ bl_int_5_150 bl_int_4_150 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c151
+ bl_int_5_151 bl_int_4_151 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c152
+ bl_int_5_152 bl_int_4_152 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c153
+ bl_int_5_153 bl_int_4_153 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c154
+ bl_int_5_154 bl_int_4_154 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c155
+ bl_int_5_155 bl_int_4_155 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c156
+ bl_int_5_156 bl_int_4_156 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c157
+ bl_int_5_157 bl_int_4_157 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c158
+ bl_int_5_158 bl_int_4_158 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c159
+ bl_int_5_159 bl_int_4_159 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c160
+ bl_int_5_160 bl_int_4_160 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c161
+ bl_int_5_161 bl_int_4_161 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c162
+ bl_int_5_162 bl_int_4_162 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c163
+ bl_int_5_163 bl_int_4_163 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c164
+ bl_int_5_164 bl_int_4_164 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c165
+ bl_int_5_165 bl_int_4_165 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c166
+ bl_int_5_166 bl_int_4_166 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c167
+ bl_int_5_167 bl_int_4_167 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c168
+ bl_int_5_168 bl_int_4_168 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c169
+ bl_int_5_169 bl_int_4_169 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c170
+ bl_int_5_170 bl_int_4_170 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c171
+ bl_int_5_171 bl_int_4_171 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c172
+ bl_int_5_172 bl_int_4_172 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c173
+ bl_int_5_173 bl_int_4_173 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c174
+ bl_int_5_174 bl_int_4_174 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c175
+ bl_int_5_175 bl_int_4_175 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c176
+ bl_int_5_176 bl_int_4_176 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c177
+ bl_int_5_177 bl_int_4_177 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c178
+ bl_int_5_178 bl_int_4_178 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c179
+ bl_int_5_179 bl_int_4_179 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c180
+ bl_int_5_180 bl_int_4_180 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c181
+ bl_int_5_181 bl_int_4_181 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c182
+ bl_int_5_182 bl_int_4_182 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r5_c183
+ bl_int_5_183 bl_int_4_183 wl_0_5 gnd
+ sram_rom_base_one_cell
Xbit_r6_c0
+ bl_int_6_0 bl_int_5_0 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c1
+ bl_int_6_1 bl_int_5_1 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c2
+ bl_int_6_2 bl_int_5_2 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c3
+ bl_int_6_3 bl_int_5_3 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c4
+ bl_int_6_4 bl_int_5_4 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c5
+ bl_int_6_5 bl_int_5_5 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c6
+ bl_int_6_6 bl_int_5_6 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c7
+ bl_int_6_7 bl_int_5_7 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c8
+ bl_int_6_8 bl_int_5_8 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c9
+ bl_int_6_9 bl_int_5_9 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c10
+ bl_int_6_10 bl_int_5_10 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c11
+ bl_int_6_11 bl_int_5_11 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c12
+ bl_int_6_12 bl_int_5_12 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c13
+ bl_int_6_13 bl_int_5_13 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c14
+ bl_int_6_14 bl_int_5_14 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c15
+ bl_int_6_15 bl_int_5_15 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c16
+ bl_int_6_16 bl_int_5_16 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c17
+ bl_int_6_17 bl_int_5_17 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c18
+ bl_int_6_18 bl_int_5_18 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c19
+ bl_int_6_19 bl_int_5_19 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c20
+ bl_int_6_20 bl_int_5_20 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c21
+ bl_int_6_21 bl_int_5_21 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c22
+ bl_int_6_22 bl_int_5_22 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c23
+ bl_int_6_23 bl_int_5_23 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c24
+ bl_int_6_24 bl_int_5_24 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c25
+ bl_int_6_25 bl_int_5_25 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c26
+ bl_int_6_26 bl_int_5_26 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c27
+ bl_int_6_27 bl_int_5_27 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c28
+ bl_int_6_28 bl_int_5_28 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c29
+ bl_int_6_29 bl_int_5_29 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c30
+ bl_int_6_30 bl_int_5_30 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c31
+ bl_int_6_31 bl_int_5_31 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c32
+ bl_int_6_32 bl_int_5_32 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c33
+ bl_int_6_33 bl_int_5_33 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c34
+ bl_int_6_34 bl_int_5_34 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c35
+ bl_int_6_35 bl_int_5_35 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c36
+ bl_int_6_36 bl_int_5_36 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c37
+ bl_int_6_37 bl_int_5_37 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c38
+ bl_int_6_38 bl_int_5_38 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c39
+ bl_int_6_39 bl_int_5_39 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c40
+ bl_int_6_40 bl_int_5_40 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c41
+ bl_int_6_41 bl_int_5_41 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c42
+ bl_int_6_42 bl_int_5_42 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c43
+ bl_int_6_43 bl_int_5_43 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c44
+ bl_int_6_44 bl_int_5_44 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c45
+ bl_int_6_45 bl_int_5_45 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c46
+ bl_int_6_46 bl_int_5_46 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c47
+ bl_int_6_47 bl_int_5_47 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c48
+ bl_int_6_48 bl_int_5_48 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c49
+ bl_int_6_49 bl_int_5_49 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c50
+ bl_int_6_50 bl_int_5_50 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c51
+ bl_int_6_51 bl_int_5_51 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c52
+ bl_int_6_52 bl_int_5_52 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c53
+ bl_int_6_53 bl_int_5_53 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c54
+ bl_int_6_54 bl_int_5_54 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c55
+ bl_int_6_55 bl_int_5_55 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c56
+ bl_int_6_56 bl_int_5_56 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c57
+ bl_int_6_57 bl_int_5_57 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c58
+ bl_int_6_58 bl_int_5_58 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c59
+ bl_int_6_59 bl_int_5_59 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c60
+ bl_int_6_60 bl_int_5_60 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c61
+ bl_int_6_61 bl_int_5_61 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c62
+ bl_int_6_62 bl_int_5_62 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c63
+ bl_int_6_63 bl_int_5_63 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c64
+ bl_int_6_64 bl_int_5_64 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c65
+ bl_int_6_65 bl_int_5_65 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c66
+ bl_int_6_66 bl_int_5_66 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c67
+ bl_int_6_67 bl_int_5_67 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c68
+ bl_int_6_68 bl_int_5_68 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c69
+ bl_int_6_69 bl_int_5_69 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c70
+ bl_int_6_70 bl_int_5_70 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c71
+ bl_int_6_71 bl_int_5_71 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c72
+ bl_int_6_72 bl_int_5_72 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c73
+ bl_int_6_73 bl_int_5_73 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c74
+ bl_int_6_74 bl_int_5_74 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c75
+ bl_int_6_75 bl_int_5_75 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c76
+ bl_int_6_76 bl_int_5_76 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c77
+ bl_int_6_77 bl_int_5_77 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c78
+ bl_int_6_78 bl_int_5_78 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c79
+ bl_int_6_79 bl_int_5_79 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c80
+ bl_int_6_80 bl_int_5_80 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c81
+ bl_int_6_81 bl_int_5_81 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c82
+ bl_int_6_82 bl_int_5_82 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c83
+ bl_int_6_83 bl_int_5_83 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c84
+ bl_int_6_84 bl_int_5_84 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c85
+ bl_int_6_85 bl_int_5_85 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c86
+ bl_int_6_86 bl_int_5_86 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c87
+ bl_int_6_87 bl_int_5_87 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c88
+ bl_int_6_88 bl_int_5_88 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c89
+ bl_int_6_89 bl_int_5_89 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c90
+ bl_int_6_90 bl_int_5_90 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c91
+ bl_int_6_91 bl_int_5_91 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c92
+ bl_int_6_92 bl_int_5_92 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c93
+ bl_int_6_93 bl_int_5_93 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c94
+ bl_int_6_94 bl_int_5_94 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c95
+ bl_int_6_95 bl_int_5_95 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c96
+ bl_int_6_96 bl_int_5_96 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c97
+ bl_int_6_97 bl_int_5_97 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c98
+ bl_int_6_98 bl_int_5_98 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c99
+ bl_int_6_99 bl_int_5_99 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c100
+ bl_int_6_100 bl_int_5_100 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c101
+ bl_int_6_101 bl_int_5_101 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c102
+ bl_int_6_102 bl_int_5_102 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c103
+ bl_int_6_103 bl_int_5_103 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c104
+ bl_int_6_104 bl_int_5_104 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c105
+ bl_int_6_105 bl_int_5_105 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c106
+ bl_int_6_106 bl_int_5_106 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c107
+ bl_int_6_107 bl_int_5_107 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c108
+ bl_int_6_108 bl_int_5_108 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c109
+ bl_int_6_109 bl_int_5_109 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c110
+ bl_int_6_110 bl_int_5_110 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c111
+ bl_int_6_111 bl_int_5_111 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c112
+ bl_int_6_112 bl_int_5_112 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c113
+ bl_int_6_113 bl_int_5_113 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c114
+ bl_int_6_114 bl_int_5_114 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c115
+ bl_int_6_115 bl_int_5_115 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c116
+ bl_int_6_116 bl_int_5_116 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c117
+ bl_int_6_117 bl_int_5_117 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c118
+ bl_int_6_118 bl_int_5_118 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c119
+ bl_int_6_119 bl_int_5_119 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c120
+ bl_int_6_120 bl_int_5_120 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c121
+ bl_int_6_121 bl_int_5_121 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c122
+ bl_int_6_122 bl_int_5_122 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c123
+ bl_int_6_123 bl_int_5_123 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c124
+ bl_int_6_124 bl_int_5_124 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c125
+ bl_int_6_125 bl_int_5_125 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c126
+ bl_int_6_126 bl_int_5_126 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c127
+ bl_int_6_127 bl_int_5_127 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c128
+ bl_int_6_128 bl_int_5_128 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c129
+ bl_int_6_129 bl_int_5_129 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c130
+ bl_int_6_130 bl_int_5_130 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c131
+ bl_int_6_131 bl_int_5_131 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c132
+ bl_int_6_132 bl_int_5_132 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c133
+ bl_int_6_133 bl_int_5_133 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c134
+ bl_int_6_134 bl_int_5_134 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c135
+ bl_int_6_135 bl_int_5_135 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c136
+ bl_int_6_136 bl_int_5_136 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c137
+ bl_int_6_137 bl_int_5_137 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c138
+ bl_int_6_138 bl_int_5_138 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c139
+ bl_int_6_139 bl_int_5_139 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c140
+ bl_int_6_140 bl_int_5_140 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c141
+ bl_int_6_141 bl_int_5_141 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c142
+ bl_int_6_142 bl_int_5_142 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c143
+ bl_int_6_143 bl_int_5_143 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c144
+ bl_int_6_144 bl_int_5_144 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c145
+ bl_int_6_145 bl_int_5_145 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c146
+ bl_int_6_146 bl_int_5_146 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c147
+ bl_int_6_147 bl_int_5_147 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c148
+ bl_int_6_148 bl_int_5_148 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c149
+ bl_int_6_149 bl_int_5_149 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c150
+ bl_int_6_150 bl_int_5_150 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c151
+ bl_int_6_151 bl_int_5_151 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c152
+ bl_int_6_152 bl_int_5_152 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c153
+ bl_int_6_153 bl_int_5_153 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c154
+ bl_int_6_154 bl_int_5_154 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c155
+ bl_int_6_155 bl_int_5_155 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c156
+ bl_int_6_156 bl_int_5_156 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c157
+ bl_int_6_157 bl_int_5_157 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c158
+ bl_int_6_158 bl_int_5_158 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c159
+ bl_int_6_159 bl_int_5_159 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c160
+ bl_int_6_160 bl_int_5_160 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c161
+ bl_int_6_161 bl_int_5_161 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c162
+ bl_int_6_162 bl_int_5_162 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c163
+ bl_int_6_163 bl_int_5_163 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c164
+ bl_int_6_164 bl_int_5_164 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c165
+ bl_int_6_165 bl_int_5_165 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c166
+ bl_int_6_166 bl_int_5_166 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c167
+ bl_int_6_167 bl_int_5_167 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c168
+ bl_int_6_168 bl_int_5_168 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c169
+ bl_int_6_169 bl_int_5_169 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c170
+ bl_int_6_170 bl_int_5_170 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c171
+ bl_int_6_171 bl_int_5_171 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c172
+ bl_int_6_172 bl_int_5_172 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c173
+ bl_int_6_173 bl_int_5_173 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c174
+ bl_int_6_174 bl_int_5_174 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c175
+ bl_int_6_175 bl_int_5_175 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c176
+ bl_int_6_176 bl_int_5_176 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c177
+ bl_int_6_177 bl_int_5_177 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c178
+ bl_int_6_178 bl_int_5_178 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c179
+ bl_int_6_179 bl_int_5_179 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c180
+ bl_int_6_180 bl_int_5_180 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c181
+ bl_int_6_181 bl_int_5_181 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c182
+ bl_int_6_182 bl_int_5_182 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r6_c183
+ bl_int_6_183 bl_int_5_183 wl_0_6 gnd
+ sram_rom_base_one_cell
Xbit_r7_c0
+ bl_int_7_0 bl_int_6_0 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c1
+ bl_int_7_1 bl_int_6_1 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c2
+ bl_int_7_2 bl_int_6_2 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c3
+ bl_int_7_3 bl_int_6_3 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c4
+ bl_int_7_4 bl_int_6_4 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c5
+ bl_int_7_5 bl_int_6_5 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c6
+ bl_int_7_6 bl_int_6_6 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c7
+ bl_int_7_7 bl_int_6_7 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c8
+ bl_int_7_8 bl_int_6_8 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c9
+ bl_int_7_9 bl_int_6_9 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c10
+ bl_int_7_10 bl_int_6_10 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c11
+ bl_int_7_11 bl_int_6_11 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c12
+ bl_int_7_12 bl_int_6_12 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c13
+ bl_int_7_13 bl_int_6_13 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c14
+ bl_int_7_14 bl_int_6_14 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c15
+ bl_int_7_15 bl_int_6_15 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c16
+ bl_int_7_16 bl_int_6_16 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c17
+ bl_int_7_17 bl_int_6_17 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c18
+ bl_int_7_18 bl_int_6_18 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c19
+ bl_int_7_19 bl_int_6_19 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c20
+ bl_int_7_20 bl_int_6_20 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c21
+ bl_int_7_21 bl_int_6_21 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c22
+ bl_int_7_22 bl_int_6_22 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c23
+ bl_int_7_23 bl_int_6_23 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c24
+ bl_int_7_24 bl_int_6_24 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c25
+ bl_int_7_25 bl_int_6_25 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c26
+ bl_int_7_26 bl_int_6_26 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c27
+ bl_int_7_27 bl_int_6_27 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c28
+ bl_int_7_28 bl_int_6_28 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c29
+ bl_int_7_29 bl_int_6_29 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c30
+ bl_int_7_30 bl_int_6_30 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c31
+ bl_int_7_31 bl_int_6_31 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c32
+ bl_int_7_32 bl_int_6_32 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c33
+ bl_int_7_33 bl_int_6_33 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c34
+ bl_int_7_34 bl_int_6_34 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c35
+ bl_int_7_35 bl_int_6_35 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c36
+ bl_int_7_36 bl_int_6_36 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c37
+ bl_int_7_37 bl_int_6_37 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c38
+ bl_int_7_38 bl_int_6_38 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c39
+ bl_int_7_39 bl_int_6_39 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c40
+ bl_int_7_40 bl_int_6_40 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c41
+ bl_int_7_41 bl_int_6_41 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c42
+ bl_int_7_42 bl_int_6_42 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c43
+ bl_int_7_43 bl_int_6_43 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c44
+ bl_int_7_44 bl_int_6_44 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c45
+ bl_int_7_45 bl_int_6_45 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c46
+ bl_int_7_46 bl_int_6_46 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c47
+ bl_int_7_47 bl_int_6_47 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c48
+ bl_int_7_48 bl_int_6_48 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c49
+ bl_int_7_49 bl_int_6_49 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c50
+ bl_int_7_50 bl_int_6_50 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c51
+ bl_int_7_51 bl_int_6_51 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c52
+ bl_int_7_52 bl_int_6_52 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c53
+ bl_int_7_53 bl_int_6_53 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c54
+ bl_int_7_54 bl_int_6_54 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c55
+ bl_int_7_55 bl_int_6_55 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c56
+ bl_int_7_56 bl_int_6_56 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c57
+ bl_int_7_57 bl_int_6_57 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c58
+ bl_int_7_58 bl_int_6_58 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c59
+ bl_int_7_59 bl_int_6_59 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c60
+ bl_int_7_60 bl_int_6_60 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c61
+ bl_int_7_61 bl_int_6_61 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c62
+ bl_int_7_62 bl_int_6_62 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c63
+ bl_int_7_63 bl_int_6_63 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c64
+ bl_int_7_64 bl_int_6_64 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c65
+ bl_int_7_65 bl_int_6_65 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c66
+ bl_int_7_66 bl_int_6_66 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c67
+ bl_int_7_67 bl_int_6_67 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c68
+ bl_int_7_68 bl_int_6_68 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c69
+ bl_int_7_69 bl_int_6_69 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c70
+ bl_int_7_70 bl_int_6_70 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c71
+ bl_int_7_71 bl_int_6_71 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c72
+ bl_int_7_72 bl_int_6_72 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c73
+ bl_int_7_73 bl_int_6_73 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c74
+ bl_int_7_74 bl_int_6_74 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c75
+ bl_int_7_75 bl_int_6_75 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c76
+ bl_int_7_76 bl_int_6_76 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c77
+ bl_int_7_77 bl_int_6_77 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c78
+ bl_int_7_78 bl_int_6_78 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c79
+ bl_int_7_79 bl_int_6_79 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c80
+ bl_int_7_80 bl_int_6_80 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c81
+ bl_int_7_81 bl_int_6_81 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c82
+ bl_int_7_82 bl_int_6_82 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c83
+ bl_int_7_83 bl_int_6_83 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c84
+ bl_int_7_84 bl_int_6_84 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c85
+ bl_int_7_85 bl_int_6_85 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c86
+ bl_int_7_86 bl_int_6_86 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c87
+ bl_int_7_87 bl_int_6_87 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c88
+ bl_int_7_88 bl_int_6_88 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c89
+ bl_int_7_89 bl_int_6_89 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c90
+ bl_int_7_90 bl_int_6_90 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c91
+ bl_int_7_91 bl_int_6_91 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c92
+ bl_int_7_92 bl_int_6_92 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c93
+ bl_int_7_93 bl_int_6_93 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c94
+ bl_int_7_94 bl_int_6_94 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c95
+ bl_int_7_95 bl_int_6_95 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c96
+ bl_int_7_96 bl_int_6_96 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c97
+ bl_int_7_97 bl_int_6_97 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c98
+ bl_int_7_98 bl_int_6_98 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c99
+ bl_int_7_99 bl_int_6_99 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c100
+ bl_int_7_100 bl_int_6_100 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c101
+ bl_int_7_101 bl_int_6_101 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c102
+ bl_int_7_102 bl_int_6_102 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c103
+ bl_int_7_103 bl_int_6_103 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c104
+ bl_int_7_104 bl_int_6_104 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c105
+ bl_int_7_105 bl_int_6_105 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c106
+ bl_int_7_106 bl_int_6_106 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c107
+ bl_int_7_107 bl_int_6_107 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c108
+ bl_int_7_108 bl_int_6_108 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c109
+ bl_int_7_109 bl_int_6_109 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c110
+ bl_int_7_110 bl_int_6_110 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c111
+ bl_int_7_111 bl_int_6_111 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c112
+ bl_int_7_112 bl_int_6_112 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c113
+ bl_int_7_113 bl_int_6_113 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c114
+ bl_int_7_114 bl_int_6_114 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c115
+ bl_int_7_115 bl_int_6_115 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c116
+ bl_int_7_116 bl_int_6_116 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c117
+ bl_int_7_117 bl_int_6_117 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c118
+ bl_int_7_118 bl_int_6_118 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c119
+ bl_int_7_119 bl_int_6_119 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c120
+ bl_int_7_120 bl_int_6_120 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c121
+ bl_int_7_121 bl_int_6_121 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c122
+ bl_int_7_122 bl_int_6_122 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c123
+ bl_int_7_123 bl_int_6_123 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c124
+ bl_int_7_124 bl_int_6_124 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c125
+ bl_int_7_125 bl_int_6_125 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c126
+ bl_int_7_126 bl_int_6_126 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c127
+ bl_int_7_127 bl_int_6_127 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c128
+ bl_int_7_128 bl_int_6_128 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c129
+ bl_int_7_129 bl_int_6_129 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c130
+ bl_int_7_130 bl_int_6_130 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c131
+ bl_int_7_131 bl_int_6_131 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c132
+ bl_int_7_132 bl_int_6_132 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c133
+ bl_int_7_133 bl_int_6_133 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c134
+ bl_int_7_134 bl_int_6_134 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c135
+ bl_int_7_135 bl_int_6_135 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c136
+ bl_int_7_136 bl_int_6_136 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c137
+ bl_int_7_137 bl_int_6_137 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c138
+ bl_int_7_138 bl_int_6_138 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c139
+ bl_int_7_139 bl_int_6_139 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c140
+ bl_int_7_140 bl_int_6_140 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c141
+ bl_int_7_141 bl_int_6_141 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c142
+ bl_int_7_142 bl_int_6_142 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c143
+ bl_int_7_143 bl_int_6_143 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c144
+ bl_int_7_144 bl_int_6_144 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c145
+ bl_int_7_145 bl_int_6_145 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c146
+ bl_int_7_146 bl_int_6_146 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c147
+ bl_int_7_147 bl_int_6_147 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c148
+ bl_int_7_148 bl_int_6_148 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c149
+ bl_int_7_149 bl_int_6_149 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c150
+ bl_int_7_150 bl_int_6_150 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c151
+ bl_int_7_151 bl_int_6_151 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c152
+ bl_int_7_152 bl_int_6_152 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c153
+ bl_int_7_153 bl_int_6_153 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c154
+ bl_int_7_154 bl_int_6_154 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c155
+ bl_int_7_155 bl_int_6_155 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c156
+ bl_int_7_156 bl_int_6_156 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c157
+ bl_int_7_157 bl_int_6_157 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c158
+ bl_int_7_158 bl_int_6_158 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c159
+ bl_int_7_159 bl_int_6_159 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c160
+ bl_int_7_160 bl_int_6_160 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c161
+ bl_int_7_161 bl_int_6_161 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c162
+ bl_int_7_162 bl_int_6_162 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c163
+ bl_int_7_163 bl_int_6_163 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c164
+ bl_int_7_164 bl_int_6_164 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c165
+ bl_int_7_165 bl_int_6_165 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c166
+ bl_int_7_166 bl_int_6_166 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c167
+ bl_int_7_167 bl_int_6_167 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c168
+ bl_int_7_168 bl_int_6_168 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c169
+ bl_int_7_169 bl_int_6_169 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c170
+ bl_int_7_170 bl_int_6_170 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c171
+ bl_int_7_171 bl_int_6_171 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c172
+ bl_int_7_172 bl_int_6_172 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c173
+ bl_int_7_173 bl_int_6_173 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c174
+ bl_int_7_174 bl_int_6_174 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c175
+ bl_int_7_175 bl_int_6_175 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c176
+ bl_int_7_176 bl_int_6_176 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c177
+ bl_int_7_177 bl_int_6_177 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c178
+ bl_int_7_178 bl_int_6_178 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c179
+ bl_int_7_179 bl_int_6_179 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c180
+ bl_int_7_180 bl_int_6_180 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c181
+ bl_int_7_181 bl_int_6_181 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c182
+ bl_int_7_182 bl_int_6_182 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r7_c183
+ bl_int_7_183 bl_int_6_183 wl_0_7 gnd
+ sram_rom_base_one_cell
Xbit_r8_c0
+ bl_int_8_0 bl_int_7_0 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c1
+ bl_int_8_1 bl_int_7_1 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c2
+ bl_int_8_2 bl_int_7_2 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c3
+ bl_int_8_3 bl_int_7_3 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c4
+ bl_int_8_4 bl_int_7_4 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c5
+ bl_int_8_5 bl_int_7_5 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c6
+ bl_int_8_6 bl_int_7_6 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c7
+ bl_int_8_7 bl_int_7_7 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c8
+ bl_int_8_8 bl_int_7_8 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c9
+ bl_int_8_9 bl_int_7_9 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c10
+ bl_int_8_10 bl_int_7_10 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c11
+ bl_int_8_11 bl_int_7_11 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c12
+ bl_int_8_12 bl_int_7_12 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c13
+ bl_int_8_13 bl_int_7_13 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c14
+ bl_int_8_14 bl_int_7_14 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c15
+ bl_int_8_15 bl_int_7_15 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c16
+ bl_int_8_16 bl_int_7_16 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c17
+ bl_int_8_17 bl_int_7_17 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c18
+ bl_int_8_18 bl_int_7_18 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c19
+ bl_int_8_19 bl_int_7_19 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c20
+ bl_int_8_20 bl_int_7_20 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c21
+ bl_int_8_21 bl_int_7_21 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c22
+ bl_int_8_22 bl_int_7_22 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c23
+ bl_int_8_23 bl_int_7_23 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c24
+ bl_int_8_24 bl_int_7_24 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c25
+ bl_int_8_25 bl_int_7_25 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c26
+ bl_int_8_26 bl_int_7_26 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c27
+ bl_int_8_27 bl_int_7_27 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c28
+ bl_int_8_28 bl_int_7_28 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c29
+ bl_int_8_29 bl_int_7_29 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c30
+ bl_int_8_30 bl_int_7_30 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c31
+ bl_int_8_31 bl_int_7_31 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c32
+ bl_int_8_32 bl_int_7_32 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c33
+ bl_int_8_33 bl_int_7_33 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c34
+ bl_int_8_34 bl_int_7_34 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c35
+ bl_int_8_35 bl_int_7_35 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c36
+ bl_int_8_36 bl_int_7_36 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c37
+ bl_int_8_37 bl_int_7_37 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c38
+ bl_int_8_38 bl_int_7_38 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c39
+ bl_int_8_39 bl_int_7_39 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c40
+ bl_int_8_40 bl_int_7_40 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c41
+ bl_int_8_41 bl_int_7_41 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c42
+ bl_int_8_42 bl_int_7_42 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c43
+ bl_int_8_43 bl_int_7_43 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c44
+ bl_int_8_44 bl_int_7_44 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c45
+ bl_int_8_45 bl_int_7_45 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c46
+ bl_int_8_46 bl_int_7_46 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c47
+ bl_int_8_47 bl_int_7_47 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c48
+ bl_int_8_48 bl_int_7_48 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c49
+ bl_int_8_49 bl_int_7_49 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c50
+ bl_int_8_50 bl_int_7_50 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c51
+ bl_int_8_51 bl_int_7_51 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c52
+ bl_int_8_52 bl_int_7_52 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c53
+ bl_int_8_53 bl_int_7_53 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c54
+ bl_int_8_54 bl_int_7_54 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c55
+ bl_int_8_55 bl_int_7_55 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c56
+ bl_int_8_56 bl_int_7_56 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c57
+ bl_int_8_57 bl_int_7_57 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c58
+ bl_int_8_58 bl_int_7_58 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c59
+ bl_int_8_59 bl_int_7_59 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c60
+ bl_int_8_60 bl_int_7_60 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c61
+ bl_int_8_61 bl_int_7_61 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c62
+ bl_int_8_62 bl_int_7_62 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c63
+ bl_int_8_63 bl_int_7_63 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c64
+ bl_int_8_64 bl_int_7_64 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c65
+ bl_int_8_65 bl_int_7_65 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c66
+ bl_int_8_66 bl_int_7_66 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c67
+ bl_int_8_67 bl_int_7_67 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c68
+ bl_int_8_68 bl_int_7_68 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c69
+ bl_int_8_69 bl_int_7_69 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c70
+ bl_int_8_70 bl_int_7_70 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c71
+ bl_int_8_71 bl_int_7_71 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c72
+ bl_int_8_72 bl_int_7_72 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c73
+ bl_int_8_73 bl_int_7_73 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c74
+ bl_int_8_74 bl_int_7_74 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c75
+ bl_int_8_75 bl_int_7_75 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c76
+ bl_int_8_76 bl_int_7_76 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c77
+ bl_int_8_77 bl_int_7_77 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c78
+ bl_int_8_78 bl_int_7_78 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c79
+ bl_int_8_79 bl_int_7_79 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c80
+ bl_int_8_80 bl_int_7_80 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c81
+ bl_int_8_81 bl_int_7_81 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c82
+ bl_int_8_82 bl_int_7_82 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c83
+ bl_int_8_83 bl_int_7_83 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c84
+ bl_int_8_84 bl_int_7_84 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c85
+ bl_int_8_85 bl_int_7_85 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c86
+ bl_int_8_86 bl_int_7_86 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c87
+ bl_int_8_87 bl_int_7_87 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c88
+ bl_int_8_88 bl_int_7_88 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c89
+ bl_int_8_89 bl_int_7_89 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c90
+ bl_int_8_90 bl_int_7_90 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c91
+ bl_int_8_91 bl_int_7_91 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c92
+ bl_int_8_92 bl_int_7_92 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c93
+ bl_int_8_93 bl_int_7_93 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c94
+ bl_int_8_94 bl_int_7_94 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c95
+ bl_int_8_95 bl_int_7_95 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c96
+ bl_int_8_96 bl_int_7_96 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c97
+ bl_int_8_97 bl_int_7_97 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c98
+ bl_int_8_98 bl_int_7_98 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c99
+ bl_int_8_99 bl_int_7_99 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c100
+ bl_int_8_100 bl_int_7_100 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c101
+ bl_int_8_101 bl_int_7_101 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c102
+ bl_int_8_102 bl_int_7_102 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c103
+ bl_int_8_103 bl_int_7_103 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c104
+ bl_int_8_104 bl_int_7_104 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c105
+ bl_int_8_105 bl_int_7_105 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c106
+ bl_int_8_106 bl_int_7_106 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c107
+ bl_int_8_107 bl_int_7_107 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c108
+ bl_int_8_108 bl_int_7_108 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c109
+ bl_int_8_109 bl_int_7_109 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c110
+ bl_int_8_110 bl_int_7_110 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c111
+ bl_int_8_111 bl_int_7_111 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c112
+ bl_int_8_112 bl_int_7_112 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c113
+ bl_int_8_113 bl_int_7_113 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c114
+ bl_int_8_114 bl_int_7_114 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c115
+ bl_int_8_115 bl_int_7_115 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c116
+ bl_int_8_116 bl_int_7_116 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c117
+ bl_int_8_117 bl_int_7_117 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c118
+ bl_int_8_118 bl_int_7_118 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c119
+ bl_int_8_119 bl_int_7_119 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c120
+ bl_int_8_120 bl_int_7_120 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c121
+ bl_int_8_121 bl_int_7_121 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c122
+ bl_int_8_122 bl_int_7_122 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c123
+ bl_int_8_123 bl_int_7_123 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c124
+ bl_int_8_124 bl_int_7_124 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c125
+ bl_int_8_125 bl_int_7_125 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c126
+ bl_int_8_126 bl_int_7_126 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c127
+ bl_int_8_127 bl_int_7_127 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c128
+ bl_int_8_128 bl_int_7_128 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c129
+ bl_int_8_129 bl_int_7_129 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c130
+ bl_int_8_130 bl_int_7_130 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c131
+ bl_int_8_131 bl_int_7_131 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c132
+ bl_int_8_132 bl_int_7_132 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c133
+ bl_int_8_133 bl_int_7_133 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c134
+ bl_int_8_134 bl_int_7_134 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c135
+ bl_int_8_135 bl_int_7_135 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c136
+ bl_int_8_136 bl_int_7_136 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c137
+ bl_int_8_137 bl_int_7_137 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c138
+ bl_int_8_138 bl_int_7_138 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c139
+ bl_int_8_139 bl_int_7_139 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c140
+ bl_int_8_140 bl_int_7_140 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c141
+ bl_int_8_141 bl_int_7_141 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c142
+ bl_int_8_142 bl_int_7_142 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c143
+ bl_int_8_143 bl_int_7_143 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c144
+ bl_int_8_144 bl_int_7_144 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c145
+ bl_int_8_145 bl_int_7_145 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c146
+ bl_int_8_146 bl_int_7_146 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c147
+ bl_int_8_147 bl_int_7_147 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c148
+ bl_int_8_148 bl_int_7_148 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c149
+ bl_int_8_149 bl_int_7_149 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c150
+ bl_int_8_150 bl_int_7_150 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c151
+ bl_int_8_151 bl_int_7_151 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c152
+ bl_int_8_152 bl_int_7_152 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c153
+ bl_int_8_153 bl_int_7_153 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c154
+ bl_int_8_154 bl_int_7_154 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c155
+ bl_int_8_155 bl_int_7_155 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c156
+ bl_int_8_156 bl_int_7_156 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c157
+ bl_int_8_157 bl_int_7_157 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c158
+ bl_int_8_158 bl_int_7_158 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c159
+ bl_int_8_159 bl_int_7_159 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c160
+ bl_int_8_160 bl_int_7_160 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c161
+ bl_int_8_161 bl_int_7_161 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c162
+ bl_int_8_162 bl_int_7_162 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c163
+ bl_int_8_163 bl_int_7_163 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c164
+ bl_int_8_164 bl_int_7_164 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c165
+ bl_int_8_165 bl_int_7_165 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c166
+ bl_int_8_166 bl_int_7_166 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c167
+ bl_int_8_167 bl_int_7_167 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c168
+ bl_int_8_168 bl_int_7_168 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c169
+ bl_int_8_169 bl_int_7_169 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c170
+ bl_int_8_170 bl_int_7_170 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c171
+ bl_int_8_171 bl_int_7_171 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c172
+ bl_int_8_172 bl_int_7_172 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c173
+ bl_int_8_173 bl_int_7_173 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c174
+ bl_int_8_174 bl_int_7_174 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c175
+ bl_int_8_175 bl_int_7_175 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c176
+ bl_int_8_176 bl_int_7_176 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c177
+ bl_int_8_177 bl_int_7_177 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c178
+ bl_int_8_178 bl_int_7_178 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c179
+ bl_int_8_179 bl_int_7_179 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c180
+ bl_int_8_180 bl_int_7_180 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c181
+ bl_int_8_181 bl_int_7_181 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c182
+ bl_int_8_182 bl_int_7_182 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r8_c183
+ bl_int_8_183 bl_int_7_183 wl_0_8 gnd
+ sram_rom_base_one_cell
Xbit_r9_c0
+ bl_int_9_0 bl_int_8_0 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c1
+ bl_int_9_1 bl_int_8_1 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c2
+ bl_int_9_2 bl_int_8_2 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c3
+ bl_int_9_3 bl_int_8_3 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c4
+ bl_int_9_4 bl_int_8_4 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c5
+ bl_int_9_5 bl_int_8_5 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c6
+ bl_int_9_6 bl_int_8_6 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c7
+ bl_int_9_7 bl_int_8_7 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c8
+ bl_int_9_8 bl_int_8_8 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c9
+ bl_int_9_9 bl_int_8_9 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c10
+ bl_int_9_10 bl_int_8_10 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c11
+ bl_int_9_11 bl_int_8_11 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c12
+ bl_int_9_12 bl_int_8_12 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c13
+ bl_int_9_13 bl_int_8_13 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c14
+ bl_int_9_14 bl_int_8_14 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c15
+ bl_int_9_15 bl_int_8_15 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c16
+ bl_int_9_16 bl_int_8_16 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c17
+ bl_int_9_17 bl_int_8_17 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c18
+ bl_int_9_18 bl_int_8_18 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c19
+ bl_int_9_19 bl_int_8_19 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c20
+ bl_int_9_20 bl_int_8_20 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c21
+ bl_int_9_21 bl_int_8_21 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c22
+ bl_int_9_22 bl_int_8_22 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c23
+ bl_int_9_23 bl_int_8_23 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c24
+ bl_int_9_24 bl_int_8_24 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c25
+ bl_int_9_25 bl_int_8_25 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c26
+ bl_int_9_26 bl_int_8_26 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c27
+ bl_int_9_27 bl_int_8_27 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c28
+ bl_int_9_28 bl_int_8_28 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c29
+ bl_int_9_29 bl_int_8_29 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c30
+ bl_int_9_30 bl_int_8_30 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c31
+ bl_int_9_31 bl_int_8_31 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c32
+ bl_int_9_32 bl_int_8_32 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c33
+ bl_int_9_33 bl_int_8_33 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c34
+ bl_int_9_34 bl_int_8_34 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c35
+ bl_int_9_35 bl_int_8_35 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c36
+ bl_int_9_36 bl_int_8_36 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c37
+ bl_int_9_37 bl_int_8_37 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c38
+ bl_int_9_38 bl_int_8_38 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c39
+ bl_int_9_39 bl_int_8_39 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c40
+ bl_int_9_40 bl_int_8_40 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c41
+ bl_int_9_41 bl_int_8_41 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c42
+ bl_int_9_42 bl_int_8_42 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c43
+ bl_int_9_43 bl_int_8_43 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c44
+ bl_int_9_44 bl_int_8_44 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c45
+ bl_int_9_45 bl_int_8_45 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c46
+ bl_int_9_46 bl_int_8_46 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c47
+ bl_int_9_47 bl_int_8_47 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c48
+ bl_int_9_48 bl_int_8_48 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c49
+ bl_int_9_49 bl_int_8_49 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c50
+ bl_int_9_50 bl_int_8_50 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c51
+ bl_int_9_51 bl_int_8_51 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c52
+ bl_int_9_52 bl_int_8_52 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c53
+ bl_int_9_53 bl_int_8_53 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c54
+ bl_int_9_54 bl_int_8_54 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c55
+ bl_int_9_55 bl_int_8_55 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c56
+ bl_int_9_56 bl_int_8_56 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c57
+ bl_int_9_57 bl_int_8_57 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c58
+ bl_int_9_58 bl_int_8_58 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c59
+ bl_int_9_59 bl_int_8_59 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c60
+ bl_int_9_60 bl_int_8_60 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c61
+ bl_int_9_61 bl_int_8_61 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c62
+ bl_int_9_62 bl_int_8_62 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c63
+ bl_int_9_63 bl_int_8_63 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c64
+ bl_int_9_64 bl_int_8_64 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c65
+ bl_int_9_65 bl_int_8_65 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c66
+ bl_int_9_66 bl_int_8_66 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c67
+ bl_int_9_67 bl_int_8_67 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c68
+ bl_int_9_68 bl_int_8_68 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c69
+ bl_int_9_69 bl_int_8_69 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c70
+ bl_int_9_70 bl_int_8_70 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c71
+ bl_int_9_71 bl_int_8_71 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c72
+ bl_int_9_72 bl_int_8_72 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c73
+ bl_int_9_73 bl_int_8_73 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c74
+ bl_int_9_74 bl_int_8_74 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c75
+ bl_int_9_75 bl_int_8_75 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c76
+ bl_int_9_76 bl_int_8_76 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c77
+ bl_int_9_77 bl_int_8_77 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c78
+ bl_int_9_78 bl_int_8_78 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c79
+ bl_int_9_79 bl_int_8_79 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c80
+ bl_int_9_80 bl_int_8_80 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c81
+ bl_int_9_81 bl_int_8_81 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c82
+ bl_int_9_82 bl_int_8_82 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c83
+ bl_int_9_83 bl_int_8_83 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c84
+ bl_int_9_84 bl_int_8_84 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c85
+ bl_int_9_85 bl_int_8_85 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c86
+ bl_int_9_86 bl_int_8_86 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c87
+ bl_int_9_87 bl_int_8_87 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c88
+ bl_int_9_88 bl_int_8_88 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c89
+ bl_int_9_89 bl_int_8_89 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c90
+ bl_int_9_90 bl_int_8_90 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c91
+ bl_int_9_91 bl_int_8_91 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c92
+ bl_int_9_92 bl_int_8_92 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c93
+ bl_int_9_93 bl_int_8_93 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c94
+ bl_int_9_94 bl_int_8_94 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c95
+ bl_int_9_95 bl_int_8_95 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c96
+ bl_int_9_96 bl_int_8_96 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c97
+ bl_int_9_97 bl_int_8_97 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c98
+ bl_int_9_98 bl_int_8_98 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c99
+ bl_int_9_99 bl_int_8_99 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c100
+ bl_int_9_100 bl_int_8_100 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c101
+ bl_int_9_101 bl_int_8_101 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c102
+ bl_int_9_102 bl_int_8_102 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c103
+ bl_int_9_103 bl_int_8_103 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c104
+ bl_int_9_104 bl_int_8_104 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c105
+ bl_int_9_105 bl_int_8_105 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c106
+ bl_int_9_106 bl_int_8_106 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c107
+ bl_int_9_107 bl_int_8_107 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c108
+ bl_int_9_108 bl_int_8_108 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c109
+ bl_int_9_109 bl_int_8_109 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c110
+ bl_int_9_110 bl_int_8_110 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c111
+ bl_int_9_111 bl_int_8_111 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c112
+ bl_int_9_112 bl_int_8_112 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c113
+ bl_int_9_113 bl_int_8_113 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c114
+ bl_int_9_114 bl_int_8_114 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c115
+ bl_int_9_115 bl_int_8_115 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c116
+ bl_int_9_116 bl_int_8_116 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c117
+ bl_int_9_117 bl_int_8_117 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c118
+ bl_int_9_118 bl_int_8_118 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c119
+ bl_int_9_119 bl_int_8_119 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c120
+ bl_int_9_120 bl_int_8_120 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c121
+ bl_int_9_121 bl_int_8_121 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c122
+ bl_int_9_122 bl_int_8_122 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c123
+ bl_int_9_123 bl_int_8_123 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c124
+ bl_int_9_124 bl_int_8_124 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c125
+ bl_int_9_125 bl_int_8_125 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c126
+ bl_int_9_126 bl_int_8_126 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c127
+ bl_int_9_127 bl_int_8_127 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c128
+ bl_int_9_128 bl_int_8_128 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c129
+ bl_int_9_129 bl_int_8_129 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c130
+ bl_int_9_130 bl_int_8_130 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c131
+ bl_int_9_131 bl_int_8_131 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c132
+ bl_int_9_132 bl_int_8_132 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c133
+ bl_int_9_133 bl_int_8_133 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c134
+ bl_int_9_134 bl_int_8_134 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c135
+ bl_int_9_135 bl_int_8_135 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c136
+ bl_int_9_136 bl_int_8_136 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c137
+ bl_int_9_137 bl_int_8_137 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c138
+ bl_int_9_138 bl_int_8_138 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c139
+ bl_int_9_139 bl_int_8_139 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c140
+ bl_int_9_140 bl_int_8_140 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c141
+ bl_int_9_141 bl_int_8_141 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c142
+ bl_int_9_142 bl_int_8_142 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c143
+ bl_int_9_143 bl_int_8_143 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c144
+ bl_int_9_144 bl_int_8_144 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c145
+ bl_int_9_145 bl_int_8_145 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c146
+ bl_int_9_146 bl_int_8_146 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c147
+ bl_int_9_147 bl_int_8_147 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c148
+ bl_int_9_148 bl_int_8_148 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c149
+ bl_int_9_149 bl_int_8_149 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c150
+ bl_int_9_150 bl_int_8_150 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c151
+ bl_int_9_151 bl_int_8_151 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c152
+ bl_int_9_152 bl_int_8_152 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c153
+ bl_int_9_153 bl_int_8_153 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c154
+ bl_int_9_154 bl_int_8_154 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c155
+ bl_int_9_155 bl_int_8_155 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c156
+ bl_int_9_156 bl_int_8_156 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c157
+ bl_int_9_157 bl_int_8_157 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c158
+ bl_int_9_158 bl_int_8_158 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c159
+ bl_int_9_159 bl_int_8_159 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c160
+ bl_int_9_160 bl_int_8_160 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c161
+ bl_int_9_161 bl_int_8_161 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c162
+ bl_int_9_162 bl_int_8_162 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c163
+ bl_int_9_163 bl_int_8_163 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c164
+ bl_int_9_164 bl_int_8_164 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c165
+ bl_int_9_165 bl_int_8_165 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c166
+ bl_int_9_166 bl_int_8_166 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c167
+ bl_int_9_167 bl_int_8_167 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c168
+ bl_int_9_168 bl_int_8_168 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c169
+ bl_int_9_169 bl_int_8_169 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c170
+ bl_int_9_170 bl_int_8_170 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c171
+ bl_int_9_171 bl_int_8_171 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c172
+ bl_int_9_172 bl_int_8_172 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c173
+ bl_int_9_173 bl_int_8_173 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c174
+ bl_int_9_174 bl_int_8_174 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c175
+ bl_int_9_175 bl_int_8_175 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c176
+ bl_int_9_176 bl_int_8_176 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c177
+ bl_int_9_177 bl_int_8_177 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c178
+ bl_int_9_178 bl_int_8_178 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c179
+ bl_int_9_179 bl_int_8_179 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c180
+ bl_int_9_180 bl_int_8_180 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c181
+ bl_int_9_181 bl_int_8_181 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c182
+ bl_int_9_182 bl_int_8_182 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r9_c183
+ bl_int_9_183 bl_int_8_183 wl_0_9 gnd
+ sram_rom_base_one_cell
Xbit_r10_c0
+ bl_int_10_0 bl_int_9_0 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c1
+ bl_int_10_1 bl_int_9_1 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c2
+ bl_int_10_2 bl_int_9_2 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c3
+ bl_int_10_3 bl_int_9_3 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c4
+ bl_int_10_4 bl_int_9_4 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c5
+ bl_int_10_5 bl_int_9_5 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c6
+ bl_int_10_6 bl_int_9_6 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c7
+ bl_int_10_7 bl_int_9_7 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c8
+ bl_int_10_8 bl_int_9_8 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c9
+ bl_int_10_9 bl_int_9_9 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c10
+ bl_int_10_10 bl_int_9_10 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c11
+ bl_int_10_11 bl_int_9_11 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c12
+ bl_int_10_12 bl_int_9_12 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c13
+ bl_int_10_13 bl_int_9_13 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c14
+ bl_int_10_14 bl_int_9_14 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c15
+ bl_int_10_15 bl_int_9_15 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c16
+ bl_int_10_16 bl_int_9_16 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c17
+ bl_int_10_17 bl_int_9_17 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c18
+ bl_int_10_18 bl_int_9_18 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c19
+ bl_int_10_19 bl_int_9_19 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c20
+ bl_int_10_20 bl_int_9_20 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c21
+ bl_int_10_21 bl_int_9_21 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c22
+ bl_int_10_22 bl_int_9_22 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c23
+ bl_int_10_23 bl_int_9_23 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c24
+ bl_int_10_24 bl_int_9_24 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c25
+ bl_int_10_25 bl_int_9_25 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c26
+ bl_int_10_26 bl_int_9_26 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c27
+ bl_int_10_27 bl_int_9_27 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c28
+ bl_int_10_28 bl_int_9_28 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c29
+ bl_int_10_29 bl_int_9_29 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c30
+ bl_int_10_30 bl_int_9_30 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c31
+ bl_int_10_31 bl_int_9_31 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c32
+ bl_int_10_32 bl_int_9_32 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c33
+ bl_int_10_33 bl_int_9_33 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c34
+ bl_int_10_34 bl_int_9_34 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c35
+ bl_int_10_35 bl_int_9_35 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c36
+ bl_int_10_36 bl_int_9_36 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c37
+ bl_int_10_37 bl_int_9_37 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c38
+ bl_int_10_38 bl_int_9_38 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c39
+ bl_int_10_39 bl_int_9_39 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c40
+ bl_int_10_40 bl_int_9_40 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c41
+ bl_int_10_41 bl_int_9_41 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c42
+ bl_int_10_42 bl_int_9_42 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c43
+ bl_int_10_43 bl_int_9_43 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c44
+ bl_int_10_44 bl_int_9_44 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c45
+ bl_int_10_45 bl_int_9_45 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c46
+ bl_int_10_46 bl_int_9_46 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c47
+ bl_int_10_47 bl_int_9_47 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c48
+ bl_int_10_48 bl_int_9_48 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c49
+ bl_int_10_49 bl_int_9_49 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c50
+ bl_int_10_50 bl_int_9_50 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c51
+ bl_int_10_51 bl_int_9_51 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c52
+ bl_int_10_52 bl_int_9_52 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c53
+ bl_int_10_53 bl_int_9_53 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c54
+ bl_int_10_54 bl_int_9_54 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c55
+ bl_int_10_55 bl_int_9_55 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c56
+ bl_int_10_56 bl_int_9_56 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c57
+ bl_int_10_57 bl_int_9_57 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c58
+ bl_int_10_58 bl_int_9_58 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c59
+ bl_int_10_59 bl_int_9_59 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c60
+ bl_int_10_60 bl_int_9_60 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c61
+ bl_int_10_61 bl_int_9_61 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c62
+ bl_int_10_62 bl_int_9_62 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c63
+ bl_int_10_63 bl_int_9_63 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c64
+ bl_int_10_64 bl_int_9_64 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c65
+ bl_int_10_65 bl_int_9_65 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c66
+ bl_int_10_66 bl_int_9_66 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c67
+ bl_int_10_67 bl_int_9_67 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c68
+ bl_int_10_68 bl_int_9_68 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c69
+ bl_int_10_69 bl_int_9_69 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c70
+ bl_int_10_70 bl_int_9_70 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c71
+ bl_int_10_71 bl_int_9_71 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c72
+ bl_int_10_72 bl_int_9_72 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c73
+ bl_int_10_73 bl_int_9_73 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c74
+ bl_int_10_74 bl_int_9_74 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c75
+ bl_int_10_75 bl_int_9_75 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c76
+ bl_int_10_76 bl_int_9_76 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c77
+ bl_int_10_77 bl_int_9_77 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c78
+ bl_int_10_78 bl_int_9_78 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c79
+ bl_int_10_79 bl_int_9_79 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c80
+ bl_int_10_80 bl_int_9_80 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c81
+ bl_int_10_81 bl_int_9_81 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c82
+ bl_int_10_82 bl_int_9_82 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c83
+ bl_int_10_83 bl_int_9_83 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c84
+ bl_int_10_84 bl_int_9_84 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c85
+ bl_int_10_85 bl_int_9_85 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c86
+ bl_int_10_86 bl_int_9_86 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c87
+ bl_int_10_87 bl_int_9_87 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c88
+ bl_int_10_88 bl_int_9_88 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c89
+ bl_int_10_89 bl_int_9_89 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c90
+ bl_int_10_90 bl_int_9_90 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c91
+ bl_int_10_91 bl_int_9_91 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c92
+ bl_int_10_92 bl_int_9_92 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c93
+ bl_int_10_93 bl_int_9_93 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c94
+ bl_int_10_94 bl_int_9_94 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c95
+ bl_int_10_95 bl_int_9_95 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c96
+ bl_int_10_96 bl_int_9_96 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c97
+ bl_int_10_97 bl_int_9_97 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c98
+ bl_int_10_98 bl_int_9_98 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c99
+ bl_int_10_99 bl_int_9_99 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c100
+ bl_int_10_100 bl_int_9_100 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c101
+ bl_int_10_101 bl_int_9_101 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c102
+ bl_int_10_102 bl_int_9_102 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c103
+ bl_int_10_103 bl_int_9_103 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c104
+ bl_int_10_104 bl_int_9_104 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c105
+ bl_int_10_105 bl_int_9_105 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c106
+ bl_int_10_106 bl_int_9_106 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c107
+ bl_int_10_107 bl_int_9_107 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c108
+ bl_int_10_108 bl_int_9_108 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c109
+ bl_int_10_109 bl_int_9_109 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c110
+ bl_int_10_110 bl_int_9_110 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c111
+ bl_int_10_111 bl_int_9_111 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c112
+ bl_int_10_112 bl_int_9_112 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c113
+ bl_int_10_113 bl_int_9_113 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c114
+ bl_int_10_114 bl_int_9_114 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c115
+ bl_int_10_115 bl_int_9_115 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c116
+ bl_int_10_116 bl_int_9_116 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c117
+ bl_int_10_117 bl_int_9_117 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c118
+ bl_int_10_118 bl_int_9_118 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c119
+ bl_int_10_119 bl_int_9_119 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c120
+ bl_int_10_120 bl_int_9_120 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c121
+ bl_int_10_121 bl_int_9_121 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c122
+ bl_int_10_122 bl_int_9_122 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c123
+ bl_int_10_123 bl_int_9_123 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c124
+ bl_int_10_124 bl_int_9_124 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c125
+ bl_int_10_125 bl_int_9_125 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c126
+ bl_int_10_126 bl_int_9_126 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c127
+ bl_int_10_127 bl_int_9_127 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c128
+ bl_int_10_128 bl_int_9_128 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c129
+ bl_int_10_129 bl_int_9_129 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c130
+ bl_int_10_130 bl_int_9_130 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c131
+ bl_int_10_131 bl_int_9_131 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c132
+ bl_int_10_132 bl_int_9_132 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c133
+ bl_int_10_133 bl_int_9_133 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c134
+ bl_int_10_134 bl_int_9_134 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c135
+ bl_int_10_135 bl_int_9_135 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c136
+ bl_int_10_136 bl_int_9_136 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c137
+ bl_int_10_137 bl_int_9_137 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c138
+ bl_int_10_138 bl_int_9_138 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c139
+ bl_int_10_139 bl_int_9_139 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c140
+ bl_int_10_140 bl_int_9_140 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c141
+ bl_int_10_141 bl_int_9_141 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c142
+ bl_int_10_142 bl_int_9_142 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c143
+ bl_int_10_143 bl_int_9_143 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c144
+ bl_int_10_144 bl_int_9_144 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c145
+ bl_int_10_145 bl_int_9_145 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c146
+ bl_int_10_146 bl_int_9_146 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c147
+ bl_int_10_147 bl_int_9_147 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c148
+ bl_int_10_148 bl_int_9_148 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c149
+ bl_int_10_149 bl_int_9_149 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c150
+ bl_int_10_150 bl_int_9_150 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c151
+ bl_int_10_151 bl_int_9_151 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c152
+ bl_int_10_152 bl_int_9_152 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c153
+ bl_int_10_153 bl_int_9_153 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c154
+ bl_int_10_154 bl_int_9_154 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c155
+ bl_int_10_155 bl_int_9_155 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c156
+ bl_int_10_156 bl_int_9_156 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c157
+ bl_int_10_157 bl_int_9_157 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c158
+ bl_int_10_158 bl_int_9_158 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c159
+ bl_int_10_159 bl_int_9_159 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c160
+ bl_int_10_160 bl_int_9_160 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c161
+ bl_int_10_161 bl_int_9_161 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c162
+ bl_int_10_162 bl_int_9_162 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c163
+ bl_int_10_163 bl_int_9_163 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c164
+ bl_int_10_164 bl_int_9_164 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c165
+ bl_int_10_165 bl_int_9_165 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c166
+ bl_int_10_166 bl_int_9_166 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c167
+ bl_int_10_167 bl_int_9_167 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c168
+ bl_int_10_168 bl_int_9_168 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c169
+ bl_int_10_169 bl_int_9_169 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c170
+ bl_int_10_170 bl_int_9_170 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c171
+ bl_int_10_171 bl_int_9_171 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c172
+ bl_int_10_172 bl_int_9_172 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c173
+ bl_int_10_173 bl_int_9_173 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c174
+ bl_int_10_174 bl_int_9_174 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c175
+ bl_int_10_175 bl_int_9_175 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c176
+ bl_int_10_176 bl_int_9_176 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c177
+ bl_int_10_177 bl_int_9_177 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c178
+ bl_int_10_178 bl_int_9_178 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c179
+ bl_int_10_179 bl_int_9_179 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c180
+ bl_int_10_180 bl_int_9_180 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c181
+ bl_int_10_181 bl_int_9_181 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c182
+ bl_int_10_182 bl_int_9_182 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r10_c183
+ bl_int_10_183 bl_int_9_183 wl_0_10 gnd
+ sram_rom_base_one_cell
Xbit_r11_c0
+ bl_int_11_0 bl_int_10_0 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c1
+ bl_int_11_1 bl_int_10_1 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c2
+ bl_int_11_2 bl_int_10_2 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c3
+ bl_int_11_3 bl_int_10_3 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c4
+ bl_int_11_4 bl_int_10_4 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c5
+ bl_int_11_5 bl_int_10_5 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c6
+ bl_int_11_6 bl_int_10_6 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c7
+ bl_int_11_7 bl_int_10_7 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c8
+ bl_int_11_8 bl_int_10_8 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c9
+ bl_int_11_9 bl_int_10_9 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c10
+ bl_int_11_10 bl_int_10_10 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c11
+ bl_int_11_11 bl_int_10_11 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c12
+ bl_int_11_12 bl_int_10_12 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c13
+ bl_int_11_13 bl_int_10_13 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c14
+ bl_int_11_14 bl_int_10_14 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c15
+ bl_int_11_15 bl_int_10_15 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c16
+ bl_int_11_16 bl_int_10_16 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c17
+ bl_int_11_17 bl_int_10_17 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c18
+ bl_int_11_18 bl_int_10_18 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c19
+ bl_int_11_19 bl_int_10_19 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c20
+ bl_int_11_20 bl_int_10_20 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c21
+ bl_int_11_21 bl_int_10_21 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c22
+ bl_int_11_22 bl_int_10_22 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c23
+ bl_int_11_23 bl_int_10_23 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c24
+ bl_int_11_24 bl_int_10_24 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c25
+ bl_int_11_25 bl_int_10_25 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c26
+ bl_int_11_26 bl_int_10_26 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c27
+ bl_int_11_27 bl_int_10_27 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c28
+ bl_int_11_28 bl_int_10_28 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c29
+ bl_int_11_29 bl_int_10_29 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c30
+ bl_int_11_30 bl_int_10_30 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c31
+ bl_int_11_31 bl_int_10_31 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c32
+ bl_int_11_32 bl_int_10_32 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c33
+ bl_int_11_33 bl_int_10_33 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c34
+ bl_int_11_34 bl_int_10_34 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c35
+ bl_int_11_35 bl_int_10_35 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c36
+ bl_int_11_36 bl_int_10_36 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c37
+ bl_int_11_37 bl_int_10_37 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c38
+ bl_int_11_38 bl_int_10_38 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c39
+ bl_int_11_39 bl_int_10_39 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c40
+ bl_int_11_40 bl_int_10_40 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c41
+ bl_int_11_41 bl_int_10_41 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c42
+ bl_int_11_42 bl_int_10_42 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c43
+ bl_int_11_43 bl_int_10_43 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c44
+ bl_int_11_44 bl_int_10_44 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c45
+ bl_int_11_45 bl_int_10_45 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c46
+ bl_int_11_46 bl_int_10_46 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c47
+ bl_int_11_47 bl_int_10_47 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c48
+ bl_int_11_48 bl_int_10_48 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c49
+ bl_int_11_49 bl_int_10_49 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c50
+ bl_int_11_50 bl_int_10_50 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c51
+ bl_int_11_51 bl_int_10_51 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c52
+ bl_int_11_52 bl_int_10_52 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c53
+ bl_int_11_53 bl_int_10_53 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c54
+ bl_int_11_54 bl_int_10_54 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c55
+ bl_int_11_55 bl_int_10_55 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c56
+ bl_int_11_56 bl_int_10_56 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c57
+ bl_int_11_57 bl_int_10_57 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c58
+ bl_int_11_58 bl_int_10_58 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c59
+ bl_int_11_59 bl_int_10_59 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c60
+ bl_int_11_60 bl_int_10_60 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c61
+ bl_int_11_61 bl_int_10_61 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c62
+ bl_int_11_62 bl_int_10_62 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c63
+ bl_int_11_63 bl_int_10_63 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c64
+ bl_int_11_64 bl_int_10_64 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c65
+ bl_int_11_65 bl_int_10_65 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c66
+ bl_int_11_66 bl_int_10_66 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c67
+ bl_int_11_67 bl_int_10_67 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c68
+ bl_int_11_68 bl_int_10_68 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c69
+ bl_int_11_69 bl_int_10_69 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c70
+ bl_int_11_70 bl_int_10_70 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c71
+ bl_int_11_71 bl_int_10_71 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c72
+ bl_int_11_72 bl_int_10_72 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c73
+ bl_int_11_73 bl_int_10_73 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c74
+ bl_int_11_74 bl_int_10_74 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c75
+ bl_int_11_75 bl_int_10_75 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c76
+ bl_int_11_76 bl_int_10_76 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c77
+ bl_int_11_77 bl_int_10_77 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c78
+ bl_int_11_78 bl_int_10_78 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c79
+ bl_int_11_79 bl_int_10_79 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c80
+ bl_int_11_80 bl_int_10_80 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c81
+ bl_int_11_81 bl_int_10_81 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c82
+ bl_int_11_82 bl_int_10_82 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c83
+ bl_int_11_83 bl_int_10_83 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c84
+ bl_int_11_84 bl_int_10_84 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c85
+ bl_int_11_85 bl_int_10_85 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c86
+ bl_int_11_86 bl_int_10_86 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c87
+ bl_int_11_87 bl_int_10_87 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c88
+ bl_int_11_88 bl_int_10_88 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c89
+ bl_int_11_89 bl_int_10_89 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c90
+ bl_int_11_90 bl_int_10_90 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c91
+ bl_int_11_91 bl_int_10_91 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c92
+ bl_int_11_92 bl_int_10_92 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c93
+ bl_int_11_93 bl_int_10_93 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c94
+ bl_int_11_94 bl_int_10_94 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c95
+ bl_int_11_95 bl_int_10_95 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c96
+ bl_int_11_96 bl_int_10_96 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c97
+ bl_int_11_97 bl_int_10_97 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c98
+ bl_int_11_98 bl_int_10_98 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c99
+ bl_int_11_99 bl_int_10_99 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c100
+ bl_int_11_100 bl_int_10_100 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c101
+ bl_int_11_101 bl_int_10_101 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c102
+ bl_int_11_102 bl_int_10_102 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c103
+ bl_int_11_103 bl_int_10_103 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c104
+ bl_int_11_104 bl_int_10_104 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c105
+ bl_int_11_105 bl_int_10_105 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c106
+ bl_int_11_106 bl_int_10_106 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c107
+ bl_int_11_107 bl_int_10_107 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c108
+ bl_int_11_108 bl_int_10_108 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c109
+ bl_int_11_109 bl_int_10_109 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c110
+ bl_int_11_110 bl_int_10_110 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c111
+ bl_int_11_111 bl_int_10_111 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c112
+ bl_int_11_112 bl_int_10_112 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c113
+ bl_int_11_113 bl_int_10_113 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c114
+ bl_int_11_114 bl_int_10_114 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c115
+ bl_int_11_115 bl_int_10_115 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c116
+ bl_int_11_116 bl_int_10_116 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c117
+ bl_int_11_117 bl_int_10_117 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c118
+ bl_int_11_118 bl_int_10_118 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c119
+ bl_int_11_119 bl_int_10_119 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c120
+ bl_int_11_120 bl_int_10_120 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c121
+ bl_int_11_121 bl_int_10_121 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c122
+ bl_int_11_122 bl_int_10_122 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c123
+ bl_int_11_123 bl_int_10_123 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c124
+ bl_int_11_124 bl_int_10_124 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c125
+ bl_int_11_125 bl_int_10_125 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c126
+ bl_int_11_126 bl_int_10_126 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c127
+ bl_int_11_127 bl_int_10_127 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c128
+ bl_int_11_128 bl_int_10_128 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c129
+ bl_int_11_129 bl_int_10_129 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c130
+ bl_int_11_130 bl_int_10_130 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c131
+ bl_int_11_131 bl_int_10_131 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c132
+ bl_int_11_132 bl_int_10_132 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c133
+ bl_int_11_133 bl_int_10_133 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c134
+ bl_int_11_134 bl_int_10_134 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c135
+ bl_int_11_135 bl_int_10_135 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c136
+ bl_int_11_136 bl_int_10_136 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c137
+ bl_int_11_137 bl_int_10_137 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c138
+ bl_int_11_138 bl_int_10_138 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c139
+ bl_int_11_139 bl_int_10_139 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c140
+ bl_int_11_140 bl_int_10_140 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c141
+ bl_int_11_141 bl_int_10_141 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c142
+ bl_int_11_142 bl_int_10_142 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c143
+ bl_int_11_143 bl_int_10_143 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c144
+ bl_int_11_144 bl_int_10_144 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c145
+ bl_int_11_145 bl_int_10_145 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c146
+ bl_int_11_146 bl_int_10_146 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c147
+ bl_int_11_147 bl_int_10_147 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c148
+ bl_int_11_148 bl_int_10_148 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c149
+ bl_int_11_149 bl_int_10_149 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c150
+ bl_int_11_150 bl_int_10_150 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c151
+ bl_int_11_151 bl_int_10_151 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c152
+ bl_int_11_152 bl_int_10_152 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c153
+ bl_int_11_153 bl_int_10_153 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c154
+ bl_int_11_154 bl_int_10_154 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c155
+ bl_int_11_155 bl_int_10_155 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c156
+ bl_int_11_156 bl_int_10_156 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c157
+ bl_int_11_157 bl_int_10_157 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c158
+ bl_int_11_158 bl_int_10_158 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c159
+ bl_int_11_159 bl_int_10_159 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c160
+ bl_int_11_160 bl_int_10_160 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c161
+ bl_int_11_161 bl_int_10_161 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c162
+ bl_int_11_162 bl_int_10_162 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c163
+ bl_int_11_163 bl_int_10_163 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c164
+ bl_int_11_164 bl_int_10_164 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c165
+ bl_int_11_165 bl_int_10_165 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c166
+ bl_int_11_166 bl_int_10_166 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c167
+ bl_int_11_167 bl_int_10_167 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c168
+ bl_int_11_168 bl_int_10_168 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c169
+ bl_int_11_169 bl_int_10_169 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c170
+ bl_int_11_170 bl_int_10_170 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c171
+ bl_int_11_171 bl_int_10_171 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c172
+ bl_int_11_172 bl_int_10_172 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c173
+ bl_int_11_173 bl_int_10_173 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c174
+ bl_int_11_174 bl_int_10_174 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c175
+ bl_int_11_175 bl_int_10_175 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c176
+ bl_int_11_176 bl_int_10_176 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c177
+ bl_int_11_177 bl_int_10_177 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c178
+ bl_int_11_178 bl_int_10_178 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c179
+ bl_int_11_179 bl_int_10_179 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c180
+ bl_int_11_180 bl_int_10_180 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c181
+ bl_int_11_181 bl_int_10_181 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c182
+ bl_int_11_182 bl_int_10_182 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r11_c183
+ bl_int_11_183 bl_int_10_183 wl_0_11 gnd
+ sram_rom_base_one_cell
Xbit_r12_c0
+ bl_int_12_0 bl_int_11_0 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c1
+ bl_int_12_1 bl_int_11_1 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c2
+ bl_int_12_2 bl_int_11_2 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c3
+ bl_int_12_3 bl_int_11_3 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c4
+ bl_int_12_4 bl_int_11_4 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c5
+ bl_int_12_5 bl_int_11_5 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c6
+ bl_int_12_6 bl_int_11_6 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c7
+ bl_int_12_7 bl_int_11_7 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c8
+ bl_int_12_8 bl_int_11_8 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c9
+ bl_int_12_9 bl_int_11_9 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c10
+ bl_int_12_10 bl_int_11_10 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c11
+ bl_int_12_11 bl_int_11_11 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c12
+ bl_int_12_12 bl_int_11_12 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c13
+ bl_int_12_13 bl_int_11_13 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c14
+ bl_int_12_14 bl_int_11_14 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c15
+ bl_int_12_15 bl_int_11_15 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c16
+ bl_int_12_16 bl_int_11_16 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c17
+ bl_int_12_17 bl_int_11_17 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c18
+ bl_int_12_18 bl_int_11_18 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c19
+ bl_int_12_19 bl_int_11_19 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c20
+ bl_int_12_20 bl_int_11_20 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c21
+ bl_int_12_21 bl_int_11_21 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c22
+ bl_int_12_22 bl_int_11_22 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c23
+ bl_int_12_23 bl_int_11_23 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c24
+ bl_int_12_24 bl_int_11_24 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c25
+ bl_int_12_25 bl_int_11_25 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c26
+ bl_int_12_26 bl_int_11_26 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c27
+ bl_int_12_27 bl_int_11_27 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c28
+ bl_int_12_28 bl_int_11_28 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c29
+ bl_int_12_29 bl_int_11_29 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c30
+ bl_int_12_30 bl_int_11_30 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c31
+ bl_int_12_31 bl_int_11_31 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c32
+ bl_int_12_32 bl_int_11_32 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c33
+ bl_int_12_33 bl_int_11_33 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c34
+ bl_int_12_34 bl_int_11_34 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c35
+ bl_int_12_35 bl_int_11_35 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c36
+ bl_int_12_36 bl_int_11_36 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c37
+ bl_int_12_37 bl_int_11_37 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c38
+ bl_int_12_38 bl_int_11_38 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c39
+ bl_int_12_39 bl_int_11_39 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c40
+ bl_int_12_40 bl_int_11_40 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c41
+ bl_int_12_41 bl_int_11_41 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c42
+ bl_int_12_42 bl_int_11_42 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c43
+ bl_int_12_43 bl_int_11_43 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c44
+ bl_int_12_44 bl_int_11_44 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c45
+ bl_int_12_45 bl_int_11_45 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c46
+ bl_int_12_46 bl_int_11_46 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c47
+ bl_int_12_47 bl_int_11_47 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c48
+ bl_int_12_48 bl_int_11_48 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c49
+ bl_int_12_49 bl_int_11_49 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c50
+ bl_int_12_50 bl_int_11_50 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c51
+ bl_int_12_51 bl_int_11_51 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c52
+ bl_int_12_52 bl_int_11_52 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c53
+ bl_int_12_53 bl_int_11_53 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c54
+ bl_int_12_54 bl_int_11_54 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c55
+ bl_int_12_55 bl_int_11_55 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c56
+ bl_int_12_56 bl_int_11_56 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c57
+ bl_int_12_57 bl_int_11_57 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c58
+ bl_int_12_58 bl_int_11_58 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c59
+ bl_int_12_59 bl_int_11_59 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c60
+ bl_int_12_60 bl_int_11_60 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c61
+ bl_int_12_61 bl_int_11_61 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c62
+ bl_int_12_62 bl_int_11_62 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c63
+ bl_int_12_63 bl_int_11_63 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c64
+ bl_int_12_64 bl_int_11_64 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c65
+ bl_int_12_65 bl_int_11_65 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c66
+ bl_int_12_66 bl_int_11_66 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c67
+ bl_int_12_67 bl_int_11_67 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c68
+ bl_int_12_68 bl_int_11_68 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c69
+ bl_int_12_69 bl_int_11_69 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c70
+ bl_int_12_70 bl_int_11_70 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c71
+ bl_int_12_71 bl_int_11_71 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c72
+ bl_int_12_72 bl_int_11_72 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c73
+ bl_int_12_73 bl_int_11_73 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c74
+ bl_int_12_74 bl_int_11_74 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c75
+ bl_int_12_75 bl_int_11_75 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c76
+ bl_int_12_76 bl_int_11_76 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c77
+ bl_int_12_77 bl_int_11_77 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c78
+ bl_int_12_78 bl_int_11_78 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c79
+ bl_int_12_79 bl_int_11_79 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c80
+ bl_int_12_80 bl_int_11_80 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c81
+ bl_int_12_81 bl_int_11_81 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c82
+ bl_int_12_82 bl_int_11_82 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c83
+ bl_int_12_83 bl_int_11_83 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c84
+ bl_int_12_84 bl_int_11_84 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c85
+ bl_int_12_85 bl_int_11_85 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c86
+ bl_int_12_86 bl_int_11_86 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c87
+ bl_int_12_87 bl_int_11_87 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c88
+ bl_int_12_88 bl_int_11_88 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c89
+ bl_int_12_89 bl_int_11_89 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c90
+ bl_int_12_90 bl_int_11_90 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c91
+ bl_int_12_91 bl_int_11_91 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c92
+ bl_int_12_92 bl_int_11_92 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c93
+ bl_int_12_93 bl_int_11_93 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c94
+ bl_int_12_94 bl_int_11_94 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c95
+ bl_int_12_95 bl_int_11_95 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c96
+ bl_int_12_96 bl_int_11_96 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c97
+ bl_int_12_97 bl_int_11_97 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c98
+ bl_int_12_98 bl_int_11_98 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c99
+ bl_int_12_99 bl_int_11_99 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c100
+ bl_int_12_100 bl_int_11_100 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c101
+ bl_int_12_101 bl_int_11_101 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c102
+ bl_int_12_102 bl_int_11_102 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c103
+ bl_int_12_103 bl_int_11_103 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c104
+ bl_int_12_104 bl_int_11_104 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c105
+ bl_int_12_105 bl_int_11_105 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c106
+ bl_int_12_106 bl_int_11_106 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c107
+ bl_int_12_107 bl_int_11_107 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c108
+ bl_int_12_108 bl_int_11_108 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c109
+ bl_int_12_109 bl_int_11_109 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c110
+ bl_int_12_110 bl_int_11_110 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c111
+ bl_int_12_111 bl_int_11_111 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c112
+ bl_int_12_112 bl_int_11_112 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c113
+ bl_int_12_113 bl_int_11_113 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c114
+ bl_int_12_114 bl_int_11_114 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c115
+ bl_int_12_115 bl_int_11_115 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c116
+ bl_int_12_116 bl_int_11_116 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c117
+ bl_int_12_117 bl_int_11_117 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c118
+ bl_int_12_118 bl_int_11_118 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c119
+ bl_int_12_119 bl_int_11_119 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c120
+ bl_int_12_120 bl_int_11_120 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c121
+ bl_int_12_121 bl_int_11_121 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c122
+ bl_int_12_122 bl_int_11_122 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c123
+ bl_int_12_123 bl_int_11_123 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c124
+ bl_int_12_124 bl_int_11_124 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c125
+ bl_int_12_125 bl_int_11_125 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c126
+ bl_int_12_126 bl_int_11_126 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c127
+ bl_int_12_127 bl_int_11_127 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c128
+ bl_int_12_128 bl_int_11_128 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c129
+ bl_int_12_129 bl_int_11_129 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c130
+ bl_int_12_130 bl_int_11_130 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c131
+ bl_int_12_131 bl_int_11_131 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c132
+ bl_int_12_132 bl_int_11_132 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c133
+ bl_int_12_133 bl_int_11_133 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c134
+ bl_int_12_134 bl_int_11_134 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c135
+ bl_int_12_135 bl_int_11_135 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c136
+ bl_int_12_136 bl_int_11_136 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c137
+ bl_int_12_137 bl_int_11_137 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c138
+ bl_int_12_138 bl_int_11_138 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c139
+ bl_int_12_139 bl_int_11_139 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c140
+ bl_int_12_140 bl_int_11_140 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c141
+ bl_int_12_141 bl_int_11_141 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c142
+ bl_int_12_142 bl_int_11_142 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c143
+ bl_int_12_143 bl_int_11_143 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c144
+ bl_int_12_144 bl_int_11_144 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c145
+ bl_int_12_145 bl_int_11_145 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c146
+ bl_int_12_146 bl_int_11_146 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c147
+ bl_int_12_147 bl_int_11_147 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c148
+ bl_int_12_148 bl_int_11_148 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c149
+ bl_int_12_149 bl_int_11_149 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c150
+ bl_int_12_150 bl_int_11_150 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c151
+ bl_int_12_151 bl_int_11_151 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c152
+ bl_int_12_152 bl_int_11_152 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c153
+ bl_int_12_153 bl_int_11_153 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c154
+ bl_int_12_154 bl_int_11_154 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c155
+ bl_int_12_155 bl_int_11_155 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c156
+ bl_int_12_156 bl_int_11_156 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c157
+ bl_int_12_157 bl_int_11_157 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c158
+ bl_int_12_158 bl_int_11_158 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c159
+ bl_int_12_159 bl_int_11_159 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c160
+ bl_int_12_160 bl_int_11_160 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c161
+ bl_int_12_161 bl_int_11_161 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c162
+ bl_int_12_162 bl_int_11_162 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c163
+ bl_int_12_163 bl_int_11_163 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c164
+ bl_int_12_164 bl_int_11_164 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c165
+ bl_int_12_165 bl_int_11_165 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c166
+ bl_int_12_166 bl_int_11_166 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c167
+ bl_int_12_167 bl_int_11_167 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c168
+ bl_int_12_168 bl_int_11_168 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c169
+ bl_int_12_169 bl_int_11_169 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c170
+ bl_int_12_170 bl_int_11_170 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c171
+ bl_int_12_171 bl_int_11_171 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c172
+ bl_int_12_172 bl_int_11_172 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c173
+ bl_int_12_173 bl_int_11_173 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c174
+ bl_int_12_174 bl_int_11_174 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c175
+ bl_int_12_175 bl_int_11_175 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c176
+ bl_int_12_176 bl_int_11_176 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c177
+ bl_int_12_177 bl_int_11_177 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c178
+ bl_int_12_178 bl_int_11_178 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c179
+ bl_int_12_179 bl_int_11_179 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c180
+ bl_int_12_180 bl_int_11_180 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c181
+ bl_int_12_181 bl_int_11_181 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c182
+ bl_int_12_182 bl_int_11_182 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r12_c183
+ bl_int_12_183 bl_int_11_183 wl_0_12 gnd
+ sram_rom_base_one_cell
Xbit_r13_c0
+ bl_int_13_0 bl_int_12_0 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c1
+ bl_int_13_1 bl_int_12_1 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c2
+ bl_int_13_2 bl_int_12_2 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c3
+ bl_int_13_3 bl_int_12_3 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c4
+ bl_int_13_4 bl_int_12_4 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c5
+ bl_int_13_5 bl_int_12_5 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c6
+ bl_int_13_6 bl_int_12_6 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c7
+ bl_int_13_7 bl_int_12_7 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c8
+ bl_int_13_8 bl_int_12_8 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c9
+ bl_int_13_9 bl_int_12_9 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c10
+ bl_int_13_10 bl_int_12_10 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c11
+ bl_int_13_11 bl_int_12_11 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c12
+ bl_int_13_12 bl_int_12_12 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c13
+ bl_int_13_13 bl_int_12_13 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c14
+ bl_int_13_14 bl_int_12_14 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c15
+ bl_int_13_15 bl_int_12_15 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c16
+ bl_int_13_16 bl_int_12_16 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c17
+ bl_int_13_17 bl_int_12_17 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c18
+ bl_int_13_18 bl_int_12_18 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c19
+ bl_int_13_19 bl_int_12_19 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c20
+ bl_int_13_20 bl_int_12_20 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c21
+ bl_int_13_21 bl_int_12_21 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c22
+ bl_int_13_22 bl_int_12_22 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c23
+ bl_int_13_23 bl_int_12_23 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c24
+ bl_int_13_24 bl_int_12_24 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c25
+ bl_int_13_25 bl_int_12_25 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c26
+ bl_int_13_26 bl_int_12_26 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c27
+ bl_int_13_27 bl_int_12_27 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c28
+ bl_int_13_28 bl_int_12_28 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c29
+ bl_int_13_29 bl_int_12_29 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c30
+ bl_int_13_30 bl_int_12_30 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c31
+ bl_int_13_31 bl_int_12_31 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c32
+ bl_int_13_32 bl_int_12_32 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c33
+ bl_int_13_33 bl_int_12_33 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c34
+ bl_int_13_34 bl_int_12_34 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c35
+ bl_int_13_35 bl_int_12_35 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c36
+ bl_int_13_36 bl_int_12_36 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c37
+ bl_int_13_37 bl_int_12_37 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c38
+ bl_int_13_38 bl_int_12_38 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c39
+ bl_int_13_39 bl_int_12_39 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c40
+ bl_int_13_40 bl_int_12_40 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c41
+ bl_int_13_41 bl_int_12_41 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c42
+ bl_int_13_42 bl_int_12_42 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c43
+ bl_int_13_43 bl_int_12_43 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c44
+ bl_int_13_44 bl_int_12_44 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c45
+ bl_int_13_45 bl_int_12_45 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c46
+ bl_int_13_46 bl_int_12_46 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c47
+ bl_int_13_47 bl_int_12_47 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c48
+ bl_int_13_48 bl_int_12_48 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c49
+ bl_int_13_49 bl_int_12_49 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c50
+ bl_int_13_50 bl_int_12_50 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c51
+ bl_int_13_51 bl_int_12_51 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c52
+ bl_int_13_52 bl_int_12_52 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c53
+ bl_int_13_53 bl_int_12_53 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c54
+ bl_int_13_54 bl_int_12_54 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c55
+ bl_int_13_55 bl_int_12_55 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c56
+ bl_int_13_56 bl_int_12_56 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c57
+ bl_int_13_57 bl_int_12_57 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c58
+ bl_int_13_58 bl_int_12_58 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c59
+ bl_int_13_59 bl_int_12_59 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c60
+ bl_int_13_60 bl_int_12_60 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c61
+ bl_int_13_61 bl_int_12_61 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c62
+ bl_int_13_62 bl_int_12_62 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c63
+ bl_int_13_63 bl_int_12_63 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c64
+ bl_int_13_64 bl_int_12_64 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c65
+ bl_int_13_65 bl_int_12_65 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c66
+ bl_int_13_66 bl_int_12_66 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c67
+ bl_int_13_67 bl_int_12_67 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c68
+ bl_int_13_68 bl_int_12_68 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c69
+ bl_int_13_69 bl_int_12_69 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c70
+ bl_int_13_70 bl_int_12_70 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c71
+ bl_int_13_71 bl_int_12_71 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c72
+ bl_int_13_72 bl_int_12_72 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c73
+ bl_int_13_73 bl_int_12_73 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c74
+ bl_int_13_74 bl_int_12_74 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c75
+ bl_int_13_75 bl_int_12_75 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c76
+ bl_int_13_76 bl_int_12_76 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c77
+ bl_int_13_77 bl_int_12_77 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c78
+ bl_int_13_78 bl_int_12_78 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c79
+ bl_int_13_79 bl_int_12_79 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c80
+ bl_int_13_80 bl_int_12_80 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c81
+ bl_int_13_81 bl_int_12_81 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c82
+ bl_int_13_82 bl_int_12_82 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c83
+ bl_int_13_83 bl_int_12_83 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c84
+ bl_int_13_84 bl_int_12_84 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c85
+ bl_int_13_85 bl_int_12_85 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c86
+ bl_int_13_86 bl_int_12_86 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c87
+ bl_int_13_87 bl_int_12_87 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c88
+ bl_int_13_88 bl_int_12_88 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c89
+ bl_int_13_89 bl_int_12_89 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c90
+ bl_int_13_90 bl_int_12_90 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c91
+ bl_int_13_91 bl_int_12_91 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c92
+ bl_int_13_92 bl_int_12_92 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c93
+ bl_int_13_93 bl_int_12_93 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c94
+ bl_int_13_94 bl_int_12_94 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c95
+ bl_int_13_95 bl_int_12_95 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c96
+ bl_int_13_96 bl_int_12_96 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c97
+ bl_int_13_97 bl_int_12_97 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c98
+ bl_int_13_98 bl_int_12_98 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c99
+ bl_int_13_99 bl_int_12_99 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c100
+ bl_int_13_100 bl_int_12_100 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c101
+ bl_int_13_101 bl_int_12_101 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c102
+ bl_int_13_102 bl_int_12_102 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c103
+ bl_int_13_103 bl_int_12_103 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c104
+ bl_int_13_104 bl_int_12_104 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c105
+ bl_int_13_105 bl_int_12_105 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c106
+ bl_int_13_106 bl_int_12_106 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c107
+ bl_int_13_107 bl_int_12_107 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c108
+ bl_int_13_108 bl_int_12_108 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c109
+ bl_int_13_109 bl_int_12_109 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c110
+ bl_int_13_110 bl_int_12_110 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c111
+ bl_int_13_111 bl_int_12_111 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c112
+ bl_int_13_112 bl_int_12_112 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c113
+ bl_int_13_113 bl_int_12_113 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c114
+ bl_int_13_114 bl_int_12_114 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c115
+ bl_int_13_115 bl_int_12_115 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c116
+ bl_int_13_116 bl_int_12_116 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c117
+ bl_int_13_117 bl_int_12_117 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c118
+ bl_int_13_118 bl_int_12_118 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c119
+ bl_int_13_119 bl_int_12_119 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c120
+ bl_int_13_120 bl_int_12_120 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c121
+ bl_int_13_121 bl_int_12_121 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c122
+ bl_int_13_122 bl_int_12_122 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c123
+ bl_int_13_123 bl_int_12_123 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c124
+ bl_int_13_124 bl_int_12_124 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c125
+ bl_int_13_125 bl_int_12_125 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c126
+ bl_int_13_126 bl_int_12_126 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c127
+ bl_int_13_127 bl_int_12_127 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c128
+ bl_int_13_128 bl_int_12_128 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c129
+ bl_int_13_129 bl_int_12_129 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c130
+ bl_int_13_130 bl_int_12_130 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c131
+ bl_int_13_131 bl_int_12_131 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c132
+ bl_int_13_132 bl_int_12_132 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c133
+ bl_int_13_133 bl_int_12_133 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c134
+ bl_int_13_134 bl_int_12_134 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c135
+ bl_int_13_135 bl_int_12_135 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c136
+ bl_int_13_136 bl_int_12_136 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c137
+ bl_int_13_137 bl_int_12_137 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c138
+ bl_int_13_138 bl_int_12_138 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c139
+ bl_int_13_139 bl_int_12_139 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c140
+ bl_int_13_140 bl_int_12_140 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c141
+ bl_int_13_141 bl_int_12_141 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c142
+ bl_int_13_142 bl_int_12_142 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c143
+ bl_int_13_143 bl_int_12_143 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c144
+ bl_int_13_144 bl_int_12_144 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c145
+ bl_int_13_145 bl_int_12_145 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c146
+ bl_int_13_146 bl_int_12_146 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c147
+ bl_int_13_147 bl_int_12_147 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c148
+ bl_int_13_148 bl_int_12_148 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c149
+ bl_int_13_149 bl_int_12_149 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c150
+ bl_int_13_150 bl_int_12_150 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c151
+ bl_int_13_151 bl_int_12_151 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c152
+ bl_int_13_152 bl_int_12_152 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c153
+ bl_int_13_153 bl_int_12_153 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c154
+ bl_int_13_154 bl_int_12_154 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c155
+ bl_int_13_155 bl_int_12_155 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c156
+ bl_int_13_156 bl_int_12_156 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c157
+ bl_int_13_157 bl_int_12_157 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c158
+ bl_int_13_158 bl_int_12_158 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c159
+ bl_int_13_159 bl_int_12_159 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c160
+ bl_int_13_160 bl_int_12_160 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c161
+ bl_int_13_161 bl_int_12_161 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c162
+ bl_int_13_162 bl_int_12_162 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c163
+ bl_int_13_163 bl_int_12_163 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c164
+ bl_int_13_164 bl_int_12_164 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c165
+ bl_int_13_165 bl_int_12_165 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c166
+ bl_int_13_166 bl_int_12_166 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c167
+ bl_int_13_167 bl_int_12_167 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c168
+ bl_int_13_168 bl_int_12_168 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c169
+ bl_int_13_169 bl_int_12_169 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c170
+ bl_int_13_170 bl_int_12_170 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c171
+ bl_int_13_171 bl_int_12_171 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c172
+ bl_int_13_172 bl_int_12_172 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c173
+ bl_int_13_173 bl_int_12_173 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c174
+ bl_int_13_174 bl_int_12_174 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c175
+ bl_int_13_175 bl_int_12_175 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c176
+ bl_int_13_176 bl_int_12_176 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c177
+ bl_int_13_177 bl_int_12_177 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c178
+ bl_int_13_178 bl_int_12_178 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c179
+ bl_int_13_179 bl_int_12_179 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c180
+ bl_int_13_180 bl_int_12_180 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c181
+ bl_int_13_181 bl_int_12_181 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c182
+ bl_int_13_182 bl_int_12_182 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r13_c183
+ bl_int_13_183 bl_int_12_183 wl_0_13 gnd
+ sram_rom_base_one_cell
Xbit_r14_c0
+ bl_int_14_0 bl_int_13_0 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c1
+ bl_int_14_1 bl_int_13_1 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c2
+ bl_int_14_2 bl_int_13_2 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c3
+ bl_int_14_3 bl_int_13_3 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c4
+ bl_int_14_4 bl_int_13_4 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c5
+ bl_int_14_5 bl_int_13_5 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c6
+ bl_int_14_6 bl_int_13_6 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c7
+ bl_int_14_7 bl_int_13_7 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c8
+ bl_int_14_8 bl_int_13_8 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c9
+ bl_int_14_9 bl_int_13_9 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c10
+ bl_int_14_10 bl_int_13_10 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c11
+ bl_int_14_11 bl_int_13_11 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c12
+ bl_int_14_12 bl_int_13_12 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c13
+ bl_int_14_13 bl_int_13_13 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c14
+ bl_int_14_14 bl_int_13_14 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c15
+ bl_int_14_15 bl_int_13_15 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c16
+ bl_int_14_16 bl_int_13_16 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c17
+ bl_int_14_17 bl_int_13_17 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c18
+ bl_int_14_18 bl_int_13_18 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c19
+ bl_int_14_19 bl_int_13_19 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c20
+ bl_int_14_20 bl_int_13_20 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c21
+ bl_int_14_21 bl_int_13_21 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c22
+ bl_int_14_22 bl_int_13_22 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c23
+ bl_int_14_23 bl_int_13_23 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c24
+ bl_int_14_24 bl_int_13_24 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c25
+ bl_int_14_25 bl_int_13_25 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c26
+ bl_int_14_26 bl_int_13_26 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c27
+ bl_int_14_27 bl_int_13_27 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c28
+ bl_int_14_28 bl_int_13_28 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c29
+ bl_int_14_29 bl_int_13_29 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c30
+ bl_int_14_30 bl_int_13_30 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c31
+ bl_int_14_31 bl_int_13_31 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c32
+ bl_int_14_32 bl_int_13_32 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c33
+ bl_int_14_33 bl_int_13_33 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c34
+ bl_int_14_34 bl_int_13_34 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c35
+ bl_int_14_35 bl_int_13_35 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c36
+ bl_int_14_36 bl_int_13_36 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c37
+ bl_int_14_37 bl_int_13_37 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c38
+ bl_int_14_38 bl_int_13_38 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c39
+ bl_int_14_39 bl_int_13_39 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c40
+ bl_int_14_40 bl_int_13_40 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c41
+ bl_int_14_41 bl_int_13_41 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c42
+ bl_int_14_42 bl_int_13_42 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c43
+ bl_int_14_43 bl_int_13_43 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c44
+ bl_int_14_44 bl_int_13_44 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c45
+ bl_int_14_45 bl_int_13_45 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c46
+ bl_int_14_46 bl_int_13_46 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c47
+ bl_int_14_47 bl_int_13_47 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c48
+ bl_int_14_48 bl_int_13_48 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c49
+ bl_int_14_49 bl_int_13_49 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c50
+ bl_int_14_50 bl_int_13_50 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c51
+ bl_int_14_51 bl_int_13_51 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c52
+ bl_int_14_52 bl_int_13_52 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c53
+ bl_int_14_53 bl_int_13_53 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c54
+ bl_int_14_54 bl_int_13_54 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c55
+ bl_int_14_55 bl_int_13_55 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c56
+ bl_int_14_56 bl_int_13_56 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c57
+ bl_int_14_57 bl_int_13_57 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c58
+ bl_int_14_58 bl_int_13_58 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c59
+ bl_int_14_59 bl_int_13_59 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c60
+ bl_int_14_60 bl_int_13_60 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c61
+ bl_int_14_61 bl_int_13_61 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c62
+ bl_int_14_62 bl_int_13_62 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c63
+ bl_int_14_63 bl_int_13_63 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c64
+ bl_int_14_64 bl_int_13_64 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c65
+ bl_int_14_65 bl_int_13_65 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c66
+ bl_int_14_66 bl_int_13_66 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c67
+ bl_int_14_67 bl_int_13_67 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c68
+ bl_int_14_68 bl_int_13_68 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c69
+ bl_int_14_69 bl_int_13_69 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c70
+ bl_int_14_70 bl_int_13_70 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c71
+ bl_int_14_71 bl_int_13_71 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c72
+ bl_int_14_72 bl_int_13_72 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c73
+ bl_int_14_73 bl_int_13_73 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c74
+ bl_int_14_74 bl_int_13_74 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c75
+ bl_int_14_75 bl_int_13_75 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c76
+ bl_int_14_76 bl_int_13_76 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c77
+ bl_int_14_77 bl_int_13_77 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c78
+ bl_int_14_78 bl_int_13_78 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c79
+ bl_int_14_79 bl_int_13_79 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c80
+ bl_int_14_80 bl_int_13_80 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c81
+ bl_int_14_81 bl_int_13_81 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c82
+ bl_int_14_82 bl_int_13_82 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c83
+ bl_int_14_83 bl_int_13_83 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c84
+ bl_int_14_84 bl_int_13_84 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c85
+ bl_int_14_85 bl_int_13_85 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c86
+ bl_int_14_86 bl_int_13_86 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c87
+ bl_int_14_87 bl_int_13_87 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c88
+ bl_int_14_88 bl_int_13_88 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c89
+ bl_int_14_89 bl_int_13_89 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c90
+ bl_int_14_90 bl_int_13_90 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c91
+ bl_int_14_91 bl_int_13_91 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c92
+ bl_int_14_92 bl_int_13_92 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c93
+ bl_int_14_93 bl_int_13_93 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c94
+ bl_int_14_94 bl_int_13_94 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c95
+ bl_int_14_95 bl_int_13_95 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c96
+ bl_int_14_96 bl_int_13_96 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c97
+ bl_int_14_97 bl_int_13_97 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c98
+ bl_int_14_98 bl_int_13_98 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c99
+ bl_int_14_99 bl_int_13_99 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c100
+ bl_int_14_100 bl_int_13_100 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c101
+ bl_int_14_101 bl_int_13_101 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c102
+ bl_int_14_102 bl_int_13_102 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c103
+ bl_int_14_103 bl_int_13_103 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c104
+ bl_int_14_104 bl_int_13_104 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c105
+ bl_int_14_105 bl_int_13_105 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c106
+ bl_int_14_106 bl_int_13_106 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c107
+ bl_int_14_107 bl_int_13_107 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c108
+ bl_int_14_108 bl_int_13_108 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c109
+ bl_int_14_109 bl_int_13_109 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c110
+ bl_int_14_110 bl_int_13_110 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c111
+ bl_int_14_111 bl_int_13_111 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c112
+ bl_int_14_112 bl_int_13_112 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c113
+ bl_int_14_113 bl_int_13_113 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c114
+ bl_int_14_114 bl_int_13_114 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c115
+ bl_int_14_115 bl_int_13_115 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c116
+ bl_int_14_116 bl_int_13_116 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c117
+ bl_int_14_117 bl_int_13_117 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c118
+ bl_int_14_118 bl_int_13_118 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c119
+ bl_int_14_119 bl_int_13_119 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c120
+ bl_int_14_120 bl_int_13_120 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c121
+ bl_int_14_121 bl_int_13_121 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c122
+ bl_int_14_122 bl_int_13_122 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c123
+ bl_int_14_123 bl_int_13_123 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c124
+ bl_int_14_124 bl_int_13_124 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c125
+ bl_int_14_125 bl_int_13_125 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c126
+ bl_int_14_126 bl_int_13_126 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c127
+ bl_int_14_127 bl_int_13_127 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c128
+ bl_int_14_128 bl_int_13_128 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c129
+ bl_int_14_129 bl_int_13_129 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c130
+ bl_int_14_130 bl_int_13_130 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c131
+ bl_int_14_131 bl_int_13_131 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c132
+ bl_int_14_132 bl_int_13_132 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c133
+ bl_int_14_133 bl_int_13_133 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c134
+ bl_int_14_134 bl_int_13_134 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c135
+ bl_int_14_135 bl_int_13_135 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c136
+ bl_int_14_136 bl_int_13_136 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c137
+ bl_int_14_137 bl_int_13_137 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c138
+ bl_int_14_138 bl_int_13_138 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c139
+ bl_int_14_139 bl_int_13_139 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c140
+ bl_int_14_140 bl_int_13_140 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c141
+ bl_int_14_141 bl_int_13_141 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c142
+ bl_int_14_142 bl_int_13_142 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c143
+ bl_int_14_143 bl_int_13_143 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c144
+ bl_int_14_144 bl_int_13_144 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c145
+ bl_int_14_145 bl_int_13_145 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c146
+ bl_int_14_146 bl_int_13_146 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c147
+ bl_int_14_147 bl_int_13_147 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c148
+ bl_int_14_148 bl_int_13_148 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c149
+ bl_int_14_149 bl_int_13_149 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c150
+ bl_int_14_150 bl_int_13_150 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c151
+ bl_int_14_151 bl_int_13_151 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c152
+ bl_int_14_152 bl_int_13_152 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c153
+ bl_int_14_153 bl_int_13_153 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c154
+ bl_int_14_154 bl_int_13_154 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c155
+ bl_int_14_155 bl_int_13_155 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c156
+ bl_int_14_156 bl_int_13_156 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c157
+ bl_int_14_157 bl_int_13_157 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c158
+ bl_int_14_158 bl_int_13_158 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c159
+ bl_int_14_159 bl_int_13_159 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c160
+ bl_int_14_160 bl_int_13_160 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c161
+ bl_int_14_161 bl_int_13_161 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c162
+ bl_int_14_162 bl_int_13_162 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c163
+ bl_int_14_163 bl_int_13_163 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c164
+ bl_int_14_164 bl_int_13_164 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c165
+ bl_int_14_165 bl_int_13_165 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c166
+ bl_int_14_166 bl_int_13_166 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c167
+ bl_int_14_167 bl_int_13_167 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c168
+ bl_int_14_168 bl_int_13_168 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c169
+ bl_int_14_169 bl_int_13_169 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c170
+ bl_int_14_170 bl_int_13_170 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c171
+ bl_int_14_171 bl_int_13_171 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c172
+ bl_int_14_172 bl_int_13_172 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c173
+ bl_int_14_173 bl_int_13_173 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c174
+ bl_int_14_174 bl_int_13_174 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c175
+ bl_int_14_175 bl_int_13_175 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c176
+ bl_int_14_176 bl_int_13_176 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c177
+ bl_int_14_177 bl_int_13_177 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c178
+ bl_int_14_178 bl_int_13_178 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c179
+ bl_int_14_179 bl_int_13_179 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c180
+ bl_int_14_180 bl_int_13_180 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c181
+ bl_int_14_181 bl_int_13_181 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c182
+ bl_int_14_182 bl_int_13_182 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r14_c183
+ bl_int_14_183 bl_int_13_183 wl_0_14 gnd
+ sram_rom_base_one_cell
Xbit_r15_c0
+ bl_int_15_0 bl_int_14_0 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c1
+ bl_int_15_1 bl_int_14_1 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c2
+ bl_int_15_2 bl_int_14_2 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c3
+ bl_int_15_3 bl_int_14_3 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c4
+ bl_int_15_4 bl_int_14_4 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c5
+ bl_int_15_5 bl_int_14_5 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c6
+ bl_int_15_6 bl_int_14_6 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c7
+ bl_int_15_7 bl_int_14_7 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c8
+ bl_int_15_8 bl_int_14_8 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c9
+ bl_int_15_9 bl_int_14_9 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c10
+ bl_int_15_10 bl_int_14_10 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c11
+ bl_int_15_11 bl_int_14_11 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c12
+ bl_int_15_12 bl_int_14_12 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c13
+ bl_int_15_13 bl_int_14_13 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c14
+ bl_int_15_14 bl_int_14_14 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c15
+ bl_int_15_15 bl_int_14_15 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c16
+ bl_int_15_16 bl_int_14_16 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c17
+ bl_int_15_17 bl_int_14_17 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c18
+ bl_int_15_18 bl_int_14_18 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c19
+ bl_int_15_19 bl_int_14_19 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c20
+ bl_int_15_20 bl_int_14_20 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c21
+ bl_int_15_21 bl_int_14_21 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c22
+ bl_int_15_22 bl_int_14_22 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c23
+ bl_int_15_23 bl_int_14_23 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c24
+ bl_int_15_24 bl_int_14_24 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c25
+ bl_int_15_25 bl_int_14_25 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c26
+ bl_int_15_26 bl_int_14_26 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c27
+ bl_int_15_27 bl_int_14_27 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c28
+ bl_int_15_28 bl_int_14_28 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c29
+ bl_int_15_29 bl_int_14_29 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c30
+ bl_int_15_30 bl_int_14_30 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c31
+ bl_int_15_31 bl_int_14_31 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c32
+ bl_int_15_32 bl_int_14_32 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c33
+ bl_int_15_33 bl_int_14_33 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c34
+ bl_int_15_34 bl_int_14_34 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c35
+ bl_int_15_35 bl_int_14_35 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c36
+ bl_int_15_36 bl_int_14_36 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c37
+ bl_int_15_37 bl_int_14_37 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c38
+ bl_int_15_38 bl_int_14_38 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c39
+ bl_int_15_39 bl_int_14_39 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c40
+ bl_int_15_40 bl_int_14_40 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c41
+ bl_int_15_41 bl_int_14_41 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c42
+ bl_int_15_42 bl_int_14_42 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c43
+ bl_int_15_43 bl_int_14_43 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c44
+ bl_int_15_44 bl_int_14_44 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c45
+ bl_int_15_45 bl_int_14_45 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c46
+ bl_int_15_46 bl_int_14_46 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c47
+ bl_int_15_47 bl_int_14_47 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c48
+ bl_int_15_48 bl_int_14_48 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c49
+ bl_int_15_49 bl_int_14_49 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c50
+ bl_int_15_50 bl_int_14_50 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c51
+ bl_int_15_51 bl_int_14_51 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c52
+ bl_int_15_52 bl_int_14_52 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c53
+ bl_int_15_53 bl_int_14_53 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c54
+ bl_int_15_54 bl_int_14_54 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c55
+ bl_int_15_55 bl_int_14_55 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c56
+ bl_int_15_56 bl_int_14_56 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c57
+ bl_int_15_57 bl_int_14_57 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c58
+ bl_int_15_58 bl_int_14_58 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c59
+ bl_int_15_59 bl_int_14_59 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c60
+ bl_int_15_60 bl_int_14_60 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c61
+ bl_int_15_61 bl_int_14_61 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c62
+ bl_int_15_62 bl_int_14_62 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c63
+ bl_int_15_63 bl_int_14_63 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c64
+ bl_int_15_64 bl_int_14_64 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c65
+ bl_int_15_65 bl_int_14_65 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c66
+ bl_int_15_66 bl_int_14_66 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c67
+ bl_int_15_67 bl_int_14_67 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c68
+ bl_int_15_68 bl_int_14_68 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c69
+ bl_int_15_69 bl_int_14_69 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c70
+ bl_int_15_70 bl_int_14_70 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c71
+ bl_int_15_71 bl_int_14_71 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c72
+ bl_int_15_72 bl_int_14_72 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c73
+ bl_int_15_73 bl_int_14_73 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c74
+ bl_int_15_74 bl_int_14_74 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c75
+ bl_int_15_75 bl_int_14_75 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c76
+ bl_int_15_76 bl_int_14_76 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c77
+ bl_int_15_77 bl_int_14_77 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c78
+ bl_int_15_78 bl_int_14_78 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c79
+ bl_int_15_79 bl_int_14_79 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c80
+ bl_int_15_80 bl_int_14_80 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c81
+ bl_int_15_81 bl_int_14_81 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c82
+ bl_int_15_82 bl_int_14_82 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c83
+ bl_int_15_83 bl_int_14_83 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c84
+ bl_int_15_84 bl_int_14_84 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c85
+ bl_int_15_85 bl_int_14_85 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c86
+ bl_int_15_86 bl_int_14_86 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c87
+ bl_int_15_87 bl_int_14_87 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c88
+ bl_int_15_88 bl_int_14_88 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c89
+ bl_int_15_89 bl_int_14_89 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c90
+ bl_int_15_90 bl_int_14_90 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c91
+ bl_int_15_91 bl_int_14_91 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c92
+ bl_int_15_92 bl_int_14_92 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c93
+ bl_int_15_93 bl_int_14_93 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c94
+ bl_int_15_94 bl_int_14_94 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c95
+ bl_int_15_95 bl_int_14_95 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c96
+ bl_int_15_96 bl_int_14_96 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c97
+ bl_int_15_97 bl_int_14_97 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c98
+ bl_int_15_98 bl_int_14_98 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c99
+ bl_int_15_99 bl_int_14_99 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c100
+ bl_int_15_100 bl_int_14_100 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c101
+ bl_int_15_101 bl_int_14_101 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c102
+ bl_int_15_102 bl_int_14_102 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c103
+ bl_int_15_103 bl_int_14_103 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c104
+ bl_int_15_104 bl_int_14_104 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c105
+ bl_int_15_105 bl_int_14_105 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c106
+ bl_int_15_106 bl_int_14_106 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c107
+ bl_int_15_107 bl_int_14_107 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c108
+ bl_int_15_108 bl_int_14_108 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c109
+ bl_int_15_109 bl_int_14_109 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c110
+ bl_int_15_110 bl_int_14_110 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c111
+ bl_int_15_111 bl_int_14_111 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c112
+ bl_int_15_112 bl_int_14_112 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c113
+ bl_int_15_113 bl_int_14_113 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c114
+ bl_int_15_114 bl_int_14_114 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c115
+ bl_int_15_115 bl_int_14_115 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c116
+ bl_int_15_116 bl_int_14_116 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c117
+ bl_int_15_117 bl_int_14_117 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c118
+ bl_int_15_118 bl_int_14_118 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c119
+ bl_int_15_119 bl_int_14_119 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c120
+ bl_int_15_120 bl_int_14_120 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c121
+ bl_int_15_121 bl_int_14_121 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c122
+ bl_int_15_122 bl_int_14_122 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c123
+ bl_int_15_123 bl_int_14_123 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c124
+ bl_int_15_124 bl_int_14_124 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c125
+ bl_int_15_125 bl_int_14_125 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c126
+ bl_int_15_126 bl_int_14_126 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c127
+ bl_int_15_127 bl_int_14_127 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c128
+ bl_int_15_128 bl_int_14_128 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c129
+ bl_int_15_129 bl_int_14_129 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c130
+ bl_int_15_130 bl_int_14_130 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c131
+ bl_int_15_131 bl_int_14_131 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c132
+ bl_int_15_132 bl_int_14_132 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c133
+ bl_int_15_133 bl_int_14_133 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c134
+ bl_int_15_134 bl_int_14_134 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c135
+ bl_int_15_135 bl_int_14_135 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c136
+ bl_int_15_136 bl_int_14_136 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c137
+ bl_int_15_137 bl_int_14_137 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c138
+ bl_int_15_138 bl_int_14_138 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c139
+ bl_int_15_139 bl_int_14_139 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c140
+ bl_int_15_140 bl_int_14_140 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c141
+ bl_int_15_141 bl_int_14_141 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c142
+ bl_int_15_142 bl_int_14_142 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c143
+ bl_int_15_143 bl_int_14_143 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c144
+ bl_int_15_144 bl_int_14_144 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c145
+ bl_int_15_145 bl_int_14_145 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c146
+ bl_int_15_146 bl_int_14_146 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c147
+ bl_int_15_147 bl_int_14_147 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c148
+ bl_int_15_148 bl_int_14_148 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c149
+ bl_int_15_149 bl_int_14_149 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c150
+ bl_int_15_150 bl_int_14_150 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c151
+ bl_int_15_151 bl_int_14_151 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c152
+ bl_int_15_152 bl_int_14_152 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c153
+ bl_int_15_153 bl_int_14_153 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c154
+ bl_int_15_154 bl_int_14_154 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c155
+ bl_int_15_155 bl_int_14_155 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c156
+ bl_int_15_156 bl_int_14_156 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c157
+ bl_int_15_157 bl_int_14_157 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c158
+ bl_int_15_158 bl_int_14_158 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c159
+ bl_int_15_159 bl_int_14_159 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c160
+ bl_int_15_160 bl_int_14_160 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c161
+ bl_int_15_161 bl_int_14_161 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c162
+ bl_int_15_162 bl_int_14_162 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c163
+ bl_int_15_163 bl_int_14_163 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c164
+ bl_int_15_164 bl_int_14_164 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c165
+ bl_int_15_165 bl_int_14_165 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c166
+ bl_int_15_166 bl_int_14_166 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c167
+ bl_int_15_167 bl_int_14_167 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c168
+ bl_int_15_168 bl_int_14_168 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c169
+ bl_int_15_169 bl_int_14_169 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c170
+ bl_int_15_170 bl_int_14_170 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c171
+ bl_int_15_171 bl_int_14_171 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c172
+ bl_int_15_172 bl_int_14_172 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c173
+ bl_int_15_173 bl_int_14_173 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c174
+ bl_int_15_174 bl_int_14_174 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c175
+ bl_int_15_175 bl_int_14_175 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c176
+ bl_int_15_176 bl_int_14_176 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c177
+ bl_int_15_177 bl_int_14_177 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c178
+ bl_int_15_178 bl_int_14_178 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c179
+ bl_int_15_179 bl_int_14_179 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c180
+ bl_int_15_180 bl_int_14_180 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c181
+ bl_int_15_181 bl_int_14_181 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c182
+ bl_int_15_182 bl_int_14_182 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r15_c183
+ bl_int_15_183 bl_int_14_183 wl_0_15 gnd
+ sram_rom_base_one_cell
Xbit_r16_c0
+ bl_int_16_0 bl_int_15_0 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c1
+ bl_int_16_1 bl_int_15_1 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c2
+ bl_int_16_2 bl_int_15_2 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c3
+ bl_int_16_3 bl_int_15_3 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c4
+ bl_int_16_4 bl_int_15_4 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c5
+ bl_int_16_5 bl_int_15_5 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c6
+ bl_int_16_6 bl_int_15_6 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c7
+ bl_int_16_7 bl_int_15_7 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c8
+ bl_int_16_8 bl_int_15_8 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c9
+ bl_int_16_9 bl_int_15_9 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c10
+ bl_int_16_10 bl_int_15_10 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c11
+ bl_int_16_11 bl_int_15_11 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c12
+ bl_int_16_12 bl_int_15_12 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c13
+ bl_int_16_13 bl_int_15_13 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c14
+ bl_int_16_14 bl_int_15_14 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c15
+ bl_int_16_15 bl_int_15_15 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c16
+ bl_int_16_16 bl_int_15_16 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c17
+ bl_int_16_17 bl_int_15_17 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c18
+ bl_int_16_18 bl_int_15_18 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c19
+ bl_int_16_19 bl_int_15_19 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c20
+ bl_int_16_20 bl_int_15_20 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c21
+ bl_int_16_21 bl_int_15_21 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c22
+ bl_int_16_22 bl_int_15_22 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c23
+ bl_int_16_23 bl_int_15_23 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c24
+ bl_int_16_24 bl_int_15_24 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c25
+ bl_int_16_25 bl_int_15_25 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c26
+ bl_int_16_26 bl_int_15_26 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c27
+ bl_int_16_27 bl_int_15_27 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c28
+ bl_int_16_28 bl_int_15_28 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c29
+ bl_int_16_29 bl_int_15_29 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c30
+ bl_int_16_30 bl_int_15_30 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c31
+ bl_int_16_31 bl_int_15_31 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c32
+ bl_int_16_32 bl_int_15_32 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c33
+ bl_int_16_33 bl_int_15_33 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c34
+ bl_int_16_34 bl_int_15_34 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c35
+ bl_int_16_35 bl_int_15_35 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c36
+ bl_int_16_36 bl_int_15_36 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c37
+ bl_int_16_37 bl_int_15_37 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c38
+ bl_int_16_38 bl_int_15_38 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c39
+ bl_int_16_39 bl_int_15_39 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c40
+ bl_int_16_40 bl_int_15_40 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c41
+ bl_int_16_41 bl_int_15_41 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c42
+ bl_int_16_42 bl_int_15_42 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c43
+ bl_int_16_43 bl_int_15_43 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c44
+ bl_int_16_44 bl_int_15_44 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c45
+ bl_int_16_45 bl_int_15_45 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c46
+ bl_int_16_46 bl_int_15_46 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c47
+ bl_int_16_47 bl_int_15_47 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c48
+ bl_int_16_48 bl_int_15_48 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c49
+ bl_int_16_49 bl_int_15_49 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c50
+ bl_int_16_50 bl_int_15_50 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c51
+ bl_int_16_51 bl_int_15_51 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c52
+ bl_int_16_52 bl_int_15_52 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c53
+ bl_int_16_53 bl_int_15_53 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c54
+ bl_int_16_54 bl_int_15_54 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c55
+ bl_int_16_55 bl_int_15_55 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c56
+ bl_int_16_56 bl_int_15_56 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c57
+ bl_int_16_57 bl_int_15_57 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c58
+ bl_int_16_58 bl_int_15_58 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c59
+ bl_int_16_59 bl_int_15_59 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c60
+ bl_int_16_60 bl_int_15_60 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c61
+ bl_int_16_61 bl_int_15_61 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c62
+ bl_int_16_62 bl_int_15_62 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c63
+ bl_int_16_63 bl_int_15_63 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c64
+ bl_int_16_64 bl_int_15_64 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c65
+ bl_int_16_65 bl_int_15_65 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c66
+ bl_int_16_66 bl_int_15_66 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c67
+ bl_int_16_67 bl_int_15_67 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c68
+ bl_int_16_68 bl_int_15_68 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c69
+ bl_int_16_69 bl_int_15_69 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c70
+ bl_int_16_70 bl_int_15_70 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c71
+ bl_int_16_71 bl_int_15_71 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c72
+ bl_int_16_72 bl_int_15_72 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c73
+ bl_int_16_73 bl_int_15_73 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c74
+ bl_int_16_74 bl_int_15_74 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c75
+ bl_int_16_75 bl_int_15_75 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c76
+ bl_int_16_76 bl_int_15_76 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c77
+ bl_int_16_77 bl_int_15_77 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c78
+ bl_int_16_78 bl_int_15_78 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c79
+ bl_int_16_79 bl_int_15_79 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c80
+ bl_int_16_80 bl_int_15_80 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c81
+ bl_int_16_81 bl_int_15_81 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c82
+ bl_int_16_82 bl_int_15_82 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c83
+ bl_int_16_83 bl_int_15_83 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c84
+ bl_int_16_84 bl_int_15_84 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c85
+ bl_int_16_85 bl_int_15_85 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c86
+ bl_int_16_86 bl_int_15_86 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c87
+ bl_int_16_87 bl_int_15_87 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c88
+ bl_int_16_88 bl_int_15_88 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c89
+ bl_int_16_89 bl_int_15_89 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c90
+ bl_int_16_90 bl_int_15_90 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c91
+ bl_int_16_91 bl_int_15_91 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c92
+ bl_int_16_92 bl_int_15_92 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c93
+ bl_int_16_93 bl_int_15_93 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c94
+ bl_int_16_94 bl_int_15_94 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c95
+ bl_int_16_95 bl_int_15_95 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c96
+ bl_int_16_96 bl_int_15_96 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c97
+ bl_int_16_97 bl_int_15_97 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c98
+ bl_int_16_98 bl_int_15_98 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c99
+ bl_int_16_99 bl_int_15_99 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c100
+ bl_int_16_100 bl_int_15_100 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c101
+ bl_int_16_101 bl_int_15_101 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c102
+ bl_int_16_102 bl_int_15_102 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c103
+ bl_int_16_103 bl_int_15_103 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c104
+ bl_int_16_104 bl_int_15_104 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c105
+ bl_int_16_105 bl_int_15_105 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c106
+ bl_int_16_106 bl_int_15_106 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c107
+ bl_int_16_107 bl_int_15_107 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c108
+ bl_int_16_108 bl_int_15_108 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c109
+ bl_int_16_109 bl_int_15_109 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c110
+ bl_int_16_110 bl_int_15_110 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c111
+ bl_int_16_111 bl_int_15_111 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c112
+ bl_int_16_112 bl_int_15_112 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c113
+ bl_int_16_113 bl_int_15_113 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c114
+ bl_int_16_114 bl_int_15_114 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c115
+ bl_int_16_115 bl_int_15_115 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c116
+ bl_int_16_116 bl_int_15_116 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c117
+ bl_int_16_117 bl_int_15_117 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c118
+ bl_int_16_118 bl_int_15_118 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c119
+ bl_int_16_119 bl_int_15_119 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c120
+ bl_int_16_120 bl_int_15_120 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c121
+ bl_int_16_121 bl_int_15_121 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c122
+ bl_int_16_122 bl_int_15_122 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c123
+ bl_int_16_123 bl_int_15_123 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c124
+ bl_int_16_124 bl_int_15_124 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c125
+ bl_int_16_125 bl_int_15_125 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c126
+ bl_int_16_126 bl_int_15_126 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c127
+ bl_int_16_127 bl_int_15_127 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c128
+ bl_int_16_128 bl_int_15_128 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c129
+ bl_int_16_129 bl_int_15_129 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c130
+ bl_int_16_130 bl_int_15_130 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c131
+ bl_int_16_131 bl_int_15_131 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c132
+ bl_int_16_132 bl_int_15_132 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c133
+ bl_int_16_133 bl_int_15_133 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c134
+ bl_int_16_134 bl_int_15_134 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c135
+ bl_int_16_135 bl_int_15_135 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c136
+ bl_int_16_136 bl_int_15_136 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c137
+ bl_int_16_137 bl_int_15_137 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c138
+ bl_int_16_138 bl_int_15_138 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c139
+ bl_int_16_139 bl_int_15_139 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c140
+ bl_int_16_140 bl_int_15_140 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c141
+ bl_int_16_141 bl_int_15_141 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c142
+ bl_int_16_142 bl_int_15_142 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c143
+ bl_int_16_143 bl_int_15_143 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c144
+ bl_int_16_144 bl_int_15_144 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c145
+ bl_int_16_145 bl_int_15_145 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c146
+ bl_int_16_146 bl_int_15_146 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c147
+ bl_int_16_147 bl_int_15_147 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c148
+ bl_int_16_148 bl_int_15_148 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c149
+ bl_int_16_149 bl_int_15_149 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c150
+ bl_int_16_150 bl_int_15_150 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c151
+ bl_int_16_151 bl_int_15_151 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c152
+ bl_int_16_152 bl_int_15_152 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c153
+ bl_int_16_153 bl_int_15_153 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c154
+ bl_int_16_154 bl_int_15_154 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c155
+ bl_int_16_155 bl_int_15_155 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c156
+ bl_int_16_156 bl_int_15_156 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c157
+ bl_int_16_157 bl_int_15_157 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c158
+ bl_int_16_158 bl_int_15_158 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c159
+ bl_int_16_159 bl_int_15_159 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c160
+ bl_int_16_160 bl_int_15_160 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c161
+ bl_int_16_161 bl_int_15_161 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c162
+ bl_int_16_162 bl_int_15_162 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c163
+ bl_int_16_163 bl_int_15_163 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c164
+ bl_int_16_164 bl_int_15_164 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c165
+ bl_int_16_165 bl_int_15_165 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c166
+ bl_int_16_166 bl_int_15_166 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c167
+ bl_int_16_167 bl_int_15_167 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c168
+ bl_int_16_168 bl_int_15_168 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c169
+ bl_int_16_169 bl_int_15_169 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c170
+ bl_int_16_170 bl_int_15_170 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c171
+ bl_int_16_171 bl_int_15_171 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c172
+ bl_int_16_172 bl_int_15_172 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c173
+ bl_int_16_173 bl_int_15_173 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c174
+ bl_int_16_174 bl_int_15_174 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c175
+ bl_int_16_175 bl_int_15_175 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c176
+ bl_int_16_176 bl_int_15_176 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c177
+ bl_int_16_177 bl_int_15_177 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c178
+ bl_int_16_178 bl_int_15_178 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c179
+ bl_int_16_179 bl_int_15_179 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c180
+ bl_int_16_180 bl_int_15_180 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c181
+ bl_int_16_181 bl_int_15_181 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c182
+ bl_int_16_182 bl_int_15_182 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r16_c183
+ bl_int_16_183 bl_int_15_183 wl_0_16 gnd
+ sram_rom_base_one_cell
Xbit_r17_c0
+ bl_int_17_0 bl_int_16_0 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c1
+ bl_int_17_1 bl_int_16_1 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c2
+ bl_int_17_2 bl_int_16_2 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c3
+ bl_int_17_3 bl_int_16_3 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c4
+ bl_int_17_4 bl_int_16_4 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c5
+ bl_int_17_5 bl_int_16_5 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c6
+ bl_int_17_6 bl_int_16_6 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c7
+ bl_int_17_7 bl_int_16_7 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c8
+ bl_int_17_8 bl_int_16_8 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c9
+ bl_int_17_9 bl_int_16_9 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c10
+ bl_int_17_10 bl_int_16_10 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c11
+ bl_int_17_11 bl_int_16_11 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c12
+ bl_int_17_12 bl_int_16_12 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c13
+ bl_int_17_13 bl_int_16_13 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c14
+ bl_int_17_14 bl_int_16_14 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c15
+ bl_int_17_15 bl_int_16_15 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c16
+ bl_int_17_16 bl_int_16_16 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c17
+ bl_int_17_17 bl_int_16_17 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c18
+ bl_int_17_18 bl_int_16_18 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c19
+ bl_int_17_19 bl_int_16_19 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c20
+ bl_int_17_20 bl_int_16_20 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c21
+ bl_int_17_21 bl_int_16_21 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c22
+ bl_int_17_22 bl_int_16_22 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c23
+ bl_int_17_23 bl_int_16_23 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c24
+ bl_int_17_24 bl_int_16_24 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c25
+ bl_int_17_25 bl_int_16_25 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c26
+ bl_int_17_26 bl_int_16_26 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c27
+ bl_int_17_27 bl_int_16_27 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c28
+ bl_int_17_28 bl_int_16_28 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c29
+ bl_int_17_29 bl_int_16_29 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c30
+ bl_int_17_30 bl_int_16_30 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c31
+ bl_int_17_31 bl_int_16_31 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c32
+ bl_int_17_32 bl_int_16_32 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c33
+ bl_int_17_33 bl_int_16_33 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c34
+ bl_int_17_34 bl_int_16_34 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c35
+ bl_int_17_35 bl_int_16_35 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c36
+ bl_int_17_36 bl_int_16_36 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c37
+ bl_int_17_37 bl_int_16_37 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c38
+ bl_int_17_38 bl_int_16_38 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c39
+ bl_int_17_39 bl_int_16_39 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c40
+ bl_int_17_40 bl_int_16_40 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c41
+ bl_int_17_41 bl_int_16_41 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c42
+ bl_int_17_42 bl_int_16_42 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c43
+ bl_int_17_43 bl_int_16_43 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c44
+ bl_int_17_44 bl_int_16_44 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c45
+ bl_int_17_45 bl_int_16_45 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c46
+ bl_int_17_46 bl_int_16_46 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c47
+ bl_int_17_47 bl_int_16_47 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c48
+ bl_int_17_48 bl_int_16_48 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c49
+ bl_int_17_49 bl_int_16_49 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c50
+ bl_int_17_50 bl_int_16_50 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c51
+ bl_int_17_51 bl_int_16_51 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c52
+ bl_int_17_52 bl_int_16_52 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c53
+ bl_int_17_53 bl_int_16_53 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c54
+ bl_int_17_54 bl_int_16_54 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c55
+ bl_int_17_55 bl_int_16_55 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c56
+ bl_int_17_56 bl_int_16_56 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c57
+ bl_int_17_57 bl_int_16_57 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c58
+ bl_int_17_58 bl_int_16_58 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c59
+ bl_int_17_59 bl_int_16_59 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c60
+ bl_int_17_60 bl_int_16_60 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c61
+ bl_int_17_61 bl_int_16_61 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c62
+ bl_int_17_62 bl_int_16_62 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c63
+ bl_int_17_63 bl_int_16_63 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c64
+ bl_int_17_64 bl_int_16_64 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c65
+ bl_int_17_65 bl_int_16_65 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c66
+ bl_int_17_66 bl_int_16_66 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c67
+ bl_int_17_67 bl_int_16_67 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c68
+ bl_int_17_68 bl_int_16_68 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c69
+ bl_int_17_69 bl_int_16_69 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c70
+ bl_int_17_70 bl_int_16_70 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c71
+ bl_int_17_71 bl_int_16_71 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c72
+ bl_int_17_72 bl_int_16_72 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c73
+ bl_int_17_73 bl_int_16_73 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c74
+ bl_int_17_74 bl_int_16_74 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c75
+ bl_int_17_75 bl_int_16_75 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c76
+ bl_int_17_76 bl_int_16_76 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c77
+ bl_int_17_77 bl_int_16_77 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c78
+ bl_int_17_78 bl_int_16_78 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c79
+ bl_int_17_79 bl_int_16_79 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c80
+ bl_int_17_80 bl_int_16_80 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c81
+ bl_int_17_81 bl_int_16_81 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c82
+ bl_int_17_82 bl_int_16_82 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c83
+ bl_int_17_83 bl_int_16_83 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c84
+ bl_int_17_84 bl_int_16_84 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c85
+ bl_int_17_85 bl_int_16_85 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c86
+ bl_int_17_86 bl_int_16_86 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c87
+ bl_int_17_87 bl_int_16_87 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c88
+ bl_int_17_88 bl_int_16_88 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c89
+ bl_int_17_89 bl_int_16_89 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c90
+ bl_int_17_90 bl_int_16_90 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c91
+ bl_int_17_91 bl_int_16_91 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c92
+ bl_int_17_92 bl_int_16_92 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c93
+ bl_int_17_93 bl_int_16_93 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c94
+ bl_int_17_94 bl_int_16_94 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c95
+ bl_int_17_95 bl_int_16_95 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c96
+ bl_int_17_96 bl_int_16_96 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c97
+ bl_int_17_97 bl_int_16_97 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c98
+ bl_int_17_98 bl_int_16_98 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c99
+ bl_int_17_99 bl_int_16_99 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c100
+ bl_int_17_100 bl_int_16_100 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c101
+ bl_int_17_101 bl_int_16_101 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c102
+ bl_int_17_102 bl_int_16_102 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c103
+ bl_int_17_103 bl_int_16_103 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c104
+ bl_int_17_104 bl_int_16_104 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c105
+ bl_int_17_105 bl_int_16_105 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c106
+ bl_int_17_106 bl_int_16_106 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c107
+ bl_int_17_107 bl_int_16_107 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c108
+ bl_int_17_108 bl_int_16_108 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c109
+ bl_int_17_109 bl_int_16_109 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c110
+ bl_int_17_110 bl_int_16_110 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c111
+ bl_int_17_111 bl_int_16_111 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c112
+ bl_int_17_112 bl_int_16_112 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c113
+ bl_int_17_113 bl_int_16_113 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c114
+ bl_int_17_114 bl_int_16_114 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c115
+ bl_int_17_115 bl_int_16_115 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c116
+ bl_int_17_116 bl_int_16_116 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c117
+ bl_int_17_117 bl_int_16_117 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c118
+ bl_int_17_118 bl_int_16_118 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c119
+ bl_int_17_119 bl_int_16_119 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c120
+ bl_int_17_120 bl_int_16_120 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c121
+ bl_int_17_121 bl_int_16_121 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c122
+ bl_int_17_122 bl_int_16_122 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c123
+ bl_int_17_123 bl_int_16_123 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c124
+ bl_int_17_124 bl_int_16_124 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c125
+ bl_int_17_125 bl_int_16_125 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c126
+ bl_int_17_126 bl_int_16_126 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c127
+ bl_int_17_127 bl_int_16_127 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c128
+ bl_int_17_128 bl_int_16_128 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c129
+ bl_int_17_129 bl_int_16_129 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c130
+ bl_int_17_130 bl_int_16_130 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c131
+ bl_int_17_131 bl_int_16_131 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c132
+ bl_int_17_132 bl_int_16_132 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c133
+ bl_int_17_133 bl_int_16_133 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c134
+ bl_int_17_134 bl_int_16_134 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c135
+ bl_int_17_135 bl_int_16_135 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c136
+ bl_int_17_136 bl_int_16_136 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c137
+ bl_int_17_137 bl_int_16_137 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c138
+ bl_int_17_138 bl_int_16_138 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c139
+ bl_int_17_139 bl_int_16_139 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c140
+ bl_int_17_140 bl_int_16_140 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c141
+ bl_int_17_141 bl_int_16_141 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c142
+ bl_int_17_142 bl_int_16_142 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c143
+ bl_int_17_143 bl_int_16_143 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c144
+ bl_int_17_144 bl_int_16_144 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c145
+ bl_int_17_145 bl_int_16_145 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c146
+ bl_int_17_146 bl_int_16_146 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c147
+ bl_int_17_147 bl_int_16_147 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c148
+ bl_int_17_148 bl_int_16_148 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c149
+ bl_int_17_149 bl_int_16_149 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c150
+ bl_int_17_150 bl_int_16_150 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c151
+ bl_int_17_151 bl_int_16_151 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c152
+ bl_int_17_152 bl_int_16_152 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c153
+ bl_int_17_153 bl_int_16_153 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c154
+ bl_int_17_154 bl_int_16_154 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c155
+ bl_int_17_155 bl_int_16_155 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c156
+ bl_int_17_156 bl_int_16_156 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c157
+ bl_int_17_157 bl_int_16_157 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c158
+ bl_int_17_158 bl_int_16_158 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c159
+ bl_int_17_159 bl_int_16_159 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c160
+ bl_int_17_160 bl_int_16_160 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c161
+ bl_int_17_161 bl_int_16_161 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c162
+ bl_int_17_162 bl_int_16_162 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c163
+ bl_int_17_163 bl_int_16_163 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c164
+ bl_int_17_164 bl_int_16_164 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c165
+ bl_int_17_165 bl_int_16_165 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c166
+ bl_int_17_166 bl_int_16_166 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c167
+ bl_int_17_167 bl_int_16_167 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c168
+ bl_int_17_168 bl_int_16_168 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c169
+ bl_int_17_169 bl_int_16_169 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c170
+ bl_int_17_170 bl_int_16_170 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c171
+ bl_int_17_171 bl_int_16_171 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c172
+ bl_int_17_172 bl_int_16_172 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c173
+ bl_int_17_173 bl_int_16_173 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c174
+ bl_int_17_174 bl_int_16_174 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c175
+ bl_int_17_175 bl_int_16_175 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c176
+ bl_int_17_176 bl_int_16_176 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c177
+ bl_int_17_177 bl_int_16_177 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c178
+ bl_int_17_178 bl_int_16_178 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c179
+ bl_int_17_179 bl_int_16_179 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c180
+ bl_int_17_180 bl_int_16_180 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c181
+ bl_int_17_181 bl_int_16_181 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c182
+ bl_int_17_182 bl_int_16_182 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r17_c183
+ bl_int_17_183 bl_int_16_183 wl_0_17 gnd
+ sram_rom_base_one_cell
Xbit_r18_c0
+ bl_int_18_0 bl_int_17_0 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c1
+ bl_int_18_1 bl_int_17_1 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c2
+ bl_int_18_2 bl_int_17_2 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c3
+ bl_int_18_3 bl_int_17_3 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c4
+ bl_int_18_4 bl_int_17_4 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c5
+ bl_int_18_5 bl_int_17_5 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c6
+ bl_int_18_6 bl_int_17_6 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c7
+ bl_int_18_7 bl_int_17_7 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c8
+ bl_int_18_8 bl_int_17_8 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c9
+ bl_int_18_9 bl_int_17_9 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c10
+ bl_int_18_10 bl_int_17_10 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c11
+ bl_int_18_11 bl_int_17_11 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c12
+ bl_int_18_12 bl_int_17_12 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c13
+ bl_int_18_13 bl_int_17_13 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c14
+ bl_int_18_14 bl_int_17_14 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c15
+ bl_int_18_15 bl_int_17_15 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c16
+ bl_int_18_16 bl_int_17_16 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c17
+ bl_int_18_17 bl_int_17_17 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c18
+ bl_int_18_18 bl_int_17_18 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c19
+ bl_int_18_19 bl_int_17_19 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c20
+ bl_int_18_20 bl_int_17_20 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c21
+ bl_int_18_21 bl_int_17_21 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c22
+ bl_int_18_22 bl_int_17_22 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c23
+ bl_int_18_23 bl_int_17_23 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c24
+ bl_int_18_24 bl_int_17_24 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c25
+ bl_int_18_25 bl_int_17_25 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c26
+ bl_int_18_26 bl_int_17_26 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c27
+ bl_int_18_27 bl_int_17_27 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c28
+ bl_int_18_28 bl_int_17_28 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c29
+ bl_int_18_29 bl_int_17_29 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c30
+ bl_int_18_30 bl_int_17_30 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c31
+ bl_int_18_31 bl_int_17_31 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c32
+ bl_int_18_32 bl_int_17_32 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c33
+ bl_int_18_33 bl_int_17_33 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c34
+ bl_int_18_34 bl_int_17_34 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c35
+ bl_int_18_35 bl_int_17_35 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c36
+ bl_int_18_36 bl_int_17_36 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c37
+ bl_int_18_37 bl_int_17_37 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c38
+ bl_int_18_38 bl_int_17_38 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c39
+ bl_int_18_39 bl_int_17_39 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c40
+ bl_int_18_40 bl_int_17_40 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c41
+ bl_int_18_41 bl_int_17_41 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c42
+ bl_int_18_42 bl_int_17_42 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c43
+ bl_int_18_43 bl_int_17_43 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c44
+ bl_int_18_44 bl_int_17_44 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c45
+ bl_int_18_45 bl_int_17_45 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c46
+ bl_int_18_46 bl_int_17_46 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c47
+ bl_int_18_47 bl_int_17_47 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c48
+ bl_int_18_48 bl_int_17_48 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c49
+ bl_int_18_49 bl_int_17_49 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c50
+ bl_int_18_50 bl_int_17_50 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c51
+ bl_int_18_51 bl_int_17_51 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c52
+ bl_int_18_52 bl_int_17_52 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c53
+ bl_int_18_53 bl_int_17_53 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c54
+ bl_int_18_54 bl_int_17_54 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c55
+ bl_int_18_55 bl_int_17_55 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c56
+ bl_int_18_56 bl_int_17_56 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c57
+ bl_int_18_57 bl_int_17_57 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c58
+ bl_int_18_58 bl_int_17_58 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c59
+ bl_int_18_59 bl_int_17_59 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c60
+ bl_int_18_60 bl_int_17_60 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c61
+ bl_int_18_61 bl_int_17_61 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c62
+ bl_int_18_62 bl_int_17_62 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c63
+ bl_int_18_63 bl_int_17_63 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c64
+ bl_int_18_64 bl_int_17_64 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c65
+ bl_int_18_65 bl_int_17_65 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c66
+ bl_int_18_66 bl_int_17_66 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c67
+ bl_int_18_67 bl_int_17_67 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c68
+ bl_int_18_68 bl_int_17_68 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c69
+ bl_int_18_69 bl_int_17_69 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c70
+ bl_int_18_70 bl_int_17_70 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c71
+ bl_int_18_71 bl_int_17_71 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c72
+ bl_int_18_72 bl_int_17_72 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c73
+ bl_int_18_73 bl_int_17_73 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c74
+ bl_int_18_74 bl_int_17_74 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c75
+ bl_int_18_75 bl_int_17_75 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c76
+ bl_int_18_76 bl_int_17_76 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c77
+ bl_int_18_77 bl_int_17_77 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c78
+ bl_int_18_78 bl_int_17_78 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c79
+ bl_int_18_79 bl_int_17_79 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c80
+ bl_int_18_80 bl_int_17_80 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c81
+ bl_int_18_81 bl_int_17_81 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c82
+ bl_int_18_82 bl_int_17_82 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c83
+ bl_int_18_83 bl_int_17_83 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c84
+ bl_int_18_84 bl_int_17_84 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c85
+ bl_int_18_85 bl_int_17_85 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c86
+ bl_int_18_86 bl_int_17_86 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c87
+ bl_int_18_87 bl_int_17_87 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c88
+ bl_int_18_88 bl_int_17_88 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c89
+ bl_int_18_89 bl_int_17_89 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c90
+ bl_int_18_90 bl_int_17_90 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c91
+ bl_int_18_91 bl_int_17_91 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c92
+ bl_int_18_92 bl_int_17_92 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c93
+ bl_int_18_93 bl_int_17_93 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c94
+ bl_int_18_94 bl_int_17_94 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c95
+ bl_int_18_95 bl_int_17_95 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c96
+ bl_int_18_96 bl_int_17_96 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c97
+ bl_int_18_97 bl_int_17_97 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c98
+ bl_int_18_98 bl_int_17_98 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c99
+ bl_int_18_99 bl_int_17_99 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c100
+ bl_int_18_100 bl_int_17_100 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c101
+ bl_int_18_101 bl_int_17_101 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c102
+ bl_int_18_102 bl_int_17_102 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c103
+ bl_int_18_103 bl_int_17_103 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c104
+ bl_int_18_104 bl_int_17_104 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c105
+ bl_int_18_105 bl_int_17_105 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c106
+ bl_int_18_106 bl_int_17_106 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c107
+ bl_int_18_107 bl_int_17_107 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c108
+ bl_int_18_108 bl_int_17_108 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c109
+ bl_int_18_109 bl_int_17_109 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c110
+ bl_int_18_110 bl_int_17_110 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c111
+ bl_int_18_111 bl_int_17_111 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c112
+ bl_int_18_112 bl_int_17_112 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c113
+ bl_int_18_113 bl_int_17_113 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c114
+ bl_int_18_114 bl_int_17_114 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c115
+ bl_int_18_115 bl_int_17_115 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c116
+ bl_int_18_116 bl_int_17_116 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c117
+ bl_int_18_117 bl_int_17_117 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c118
+ bl_int_18_118 bl_int_17_118 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c119
+ bl_int_18_119 bl_int_17_119 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c120
+ bl_int_18_120 bl_int_17_120 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c121
+ bl_int_18_121 bl_int_17_121 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c122
+ bl_int_18_122 bl_int_17_122 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c123
+ bl_int_18_123 bl_int_17_123 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c124
+ bl_int_18_124 bl_int_17_124 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c125
+ bl_int_18_125 bl_int_17_125 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c126
+ bl_int_18_126 bl_int_17_126 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c127
+ bl_int_18_127 bl_int_17_127 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c128
+ bl_int_18_128 bl_int_17_128 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c129
+ bl_int_18_129 bl_int_17_129 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c130
+ bl_int_18_130 bl_int_17_130 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c131
+ bl_int_18_131 bl_int_17_131 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c132
+ bl_int_18_132 bl_int_17_132 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c133
+ bl_int_18_133 bl_int_17_133 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c134
+ bl_int_18_134 bl_int_17_134 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c135
+ bl_int_18_135 bl_int_17_135 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c136
+ bl_int_18_136 bl_int_17_136 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c137
+ bl_int_18_137 bl_int_17_137 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c138
+ bl_int_18_138 bl_int_17_138 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c139
+ bl_int_18_139 bl_int_17_139 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c140
+ bl_int_18_140 bl_int_17_140 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c141
+ bl_int_18_141 bl_int_17_141 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c142
+ bl_int_18_142 bl_int_17_142 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c143
+ bl_int_18_143 bl_int_17_143 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c144
+ bl_int_18_144 bl_int_17_144 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c145
+ bl_int_18_145 bl_int_17_145 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c146
+ bl_int_18_146 bl_int_17_146 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c147
+ bl_int_18_147 bl_int_17_147 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c148
+ bl_int_18_148 bl_int_17_148 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c149
+ bl_int_18_149 bl_int_17_149 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c150
+ bl_int_18_150 bl_int_17_150 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c151
+ bl_int_18_151 bl_int_17_151 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c152
+ bl_int_18_152 bl_int_17_152 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c153
+ bl_int_18_153 bl_int_17_153 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c154
+ bl_int_18_154 bl_int_17_154 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c155
+ bl_int_18_155 bl_int_17_155 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c156
+ bl_int_18_156 bl_int_17_156 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c157
+ bl_int_18_157 bl_int_17_157 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c158
+ bl_int_18_158 bl_int_17_158 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c159
+ bl_int_18_159 bl_int_17_159 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c160
+ bl_int_18_160 bl_int_17_160 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c161
+ bl_int_18_161 bl_int_17_161 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c162
+ bl_int_18_162 bl_int_17_162 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c163
+ bl_int_18_163 bl_int_17_163 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c164
+ bl_int_18_164 bl_int_17_164 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c165
+ bl_int_18_165 bl_int_17_165 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c166
+ bl_int_18_166 bl_int_17_166 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c167
+ bl_int_18_167 bl_int_17_167 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c168
+ bl_int_18_168 bl_int_17_168 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c169
+ bl_int_18_169 bl_int_17_169 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c170
+ bl_int_18_170 bl_int_17_170 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c171
+ bl_int_18_171 bl_int_17_171 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c172
+ bl_int_18_172 bl_int_17_172 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c173
+ bl_int_18_173 bl_int_17_173 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c174
+ bl_int_18_174 bl_int_17_174 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c175
+ bl_int_18_175 bl_int_17_175 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c176
+ bl_int_18_176 bl_int_17_176 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c177
+ bl_int_18_177 bl_int_17_177 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c178
+ bl_int_18_178 bl_int_17_178 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c179
+ bl_int_18_179 bl_int_17_179 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c180
+ bl_int_18_180 bl_int_17_180 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c181
+ bl_int_18_181 bl_int_17_181 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c182
+ bl_int_18_182 bl_int_17_182 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r18_c183
+ bl_int_18_183 bl_int_17_183 wl_0_18 gnd
+ sram_rom_base_one_cell
Xbit_r19_c0
+ bl_int_19_0 bl_int_18_0 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c1
+ bl_int_19_1 bl_int_18_1 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c2
+ bl_int_19_2 bl_int_18_2 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c3
+ bl_int_19_3 bl_int_18_3 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c4
+ bl_int_19_4 bl_int_18_4 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c5
+ bl_int_19_5 bl_int_18_5 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c6
+ bl_int_19_6 bl_int_18_6 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c7
+ bl_int_19_7 bl_int_18_7 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c8
+ bl_int_19_8 bl_int_18_8 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c9
+ bl_int_19_9 bl_int_18_9 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c10
+ bl_int_19_10 bl_int_18_10 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c11
+ bl_int_19_11 bl_int_18_11 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c12
+ bl_int_19_12 bl_int_18_12 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c13
+ bl_int_19_13 bl_int_18_13 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c14
+ bl_int_19_14 bl_int_18_14 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c15
+ bl_int_19_15 bl_int_18_15 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c16
+ bl_int_19_16 bl_int_18_16 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c17
+ bl_int_19_17 bl_int_18_17 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c18
+ bl_int_19_18 bl_int_18_18 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c19
+ bl_int_19_19 bl_int_18_19 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c20
+ bl_int_19_20 bl_int_18_20 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c21
+ bl_int_19_21 bl_int_18_21 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c22
+ bl_int_19_22 bl_int_18_22 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c23
+ bl_int_19_23 bl_int_18_23 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c24
+ bl_int_19_24 bl_int_18_24 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c25
+ bl_int_19_25 bl_int_18_25 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c26
+ bl_int_19_26 bl_int_18_26 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c27
+ bl_int_19_27 bl_int_18_27 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c28
+ bl_int_19_28 bl_int_18_28 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c29
+ bl_int_19_29 bl_int_18_29 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c30
+ bl_int_19_30 bl_int_18_30 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c31
+ bl_int_19_31 bl_int_18_31 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c32
+ bl_int_19_32 bl_int_18_32 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c33
+ bl_int_19_33 bl_int_18_33 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c34
+ bl_int_19_34 bl_int_18_34 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c35
+ bl_int_19_35 bl_int_18_35 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c36
+ bl_int_19_36 bl_int_18_36 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c37
+ bl_int_19_37 bl_int_18_37 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c38
+ bl_int_19_38 bl_int_18_38 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c39
+ bl_int_19_39 bl_int_18_39 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c40
+ bl_int_19_40 bl_int_18_40 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c41
+ bl_int_19_41 bl_int_18_41 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c42
+ bl_int_19_42 bl_int_18_42 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c43
+ bl_int_19_43 bl_int_18_43 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c44
+ bl_int_19_44 bl_int_18_44 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c45
+ bl_int_19_45 bl_int_18_45 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c46
+ bl_int_19_46 bl_int_18_46 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c47
+ bl_int_19_47 bl_int_18_47 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c48
+ bl_int_19_48 bl_int_18_48 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c49
+ bl_int_19_49 bl_int_18_49 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c50
+ bl_int_19_50 bl_int_18_50 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c51
+ bl_int_19_51 bl_int_18_51 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c52
+ bl_int_19_52 bl_int_18_52 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c53
+ bl_int_19_53 bl_int_18_53 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c54
+ bl_int_19_54 bl_int_18_54 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c55
+ bl_int_19_55 bl_int_18_55 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c56
+ bl_int_19_56 bl_int_18_56 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c57
+ bl_int_19_57 bl_int_18_57 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c58
+ bl_int_19_58 bl_int_18_58 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c59
+ bl_int_19_59 bl_int_18_59 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c60
+ bl_int_19_60 bl_int_18_60 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c61
+ bl_int_19_61 bl_int_18_61 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c62
+ bl_int_19_62 bl_int_18_62 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c63
+ bl_int_19_63 bl_int_18_63 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c64
+ bl_int_19_64 bl_int_18_64 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c65
+ bl_int_19_65 bl_int_18_65 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c66
+ bl_int_19_66 bl_int_18_66 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c67
+ bl_int_19_67 bl_int_18_67 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c68
+ bl_int_19_68 bl_int_18_68 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c69
+ bl_int_19_69 bl_int_18_69 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c70
+ bl_int_19_70 bl_int_18_70 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c71
+ bl_int_19_71 bl_int_18_71 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c72
+ bl_int_19_72 bl_int_18_72 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c73
+ bl_int_19_73 bl_int_18_73 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c74
+ bl_int_19_74 bl_int_18_74 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c75
+ bl_int_19_75 bl_int_18_75 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c76
+ bl_int_19_76 bl_int_18_76 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c77
+ bl_int_19_77 bl_int_18_77 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c78
+ bl_int_19_78 bl_int_18_78 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c79
+ bl_int_19_79 bl_int_18_79 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c80
+ bl_int_19_80 bl_int_18_80 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c81
+ bl_int_19_81 bl_int_18_81 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c82
+ bl_int_19_82 bl_int_18_82 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c83
+ bl_int_19_83 bl_int_18_83 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c84
+ bl_int_19_84 bl_int_18_84 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c85
+ bl_int_19_85 bl_int_18_85 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c86
+ bl_int_19_86 bl_int_18_86 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c87
+ bl_int_19_87 bl_int_18_87 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c88
+ bl_int_19_88 bl_int_18_88 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c89
+ bl_int_19_89 bl_int_18_89 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c90
+ bl_int_19_90 bl_int_18_90 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c91
+ bl_int_19_91 bl_int_18_91 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c92
+ bl_int_19_92 bl_int_18_92 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c93
+ bl_int_19_93 bl_int_18_93 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c94
+ bl_int_19_94 bl_int_18_94 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c95
+ bl_int_19_95 bl_int_18_95 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c96
+ bl_int_19_96 bl_int_18_96 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c97
+ bl_int_19_97 bl_int_18_97 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c98
+ bl_int_19_98 bl_int_18_98 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c99
+ bl_int_19_99 bl_int_18_99 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c100
+ bl_int_19_100 bl_int_18_100 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c101
+ bl_int_19_101 bl_int_18_101 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c102
+ bl_int_19_102 bl_int_18_102 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c103
+ bl_int_19_103 bl_int_18_103 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c104
+ bl_int_19_104 bl_int_18_104 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c105
+ bl_int_19_105 bl_int_18_105 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c106
+ bl_int_19_106 bl_int_18_106 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c107
+ bl_int_19_107 bl_int_18_107 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c108
+ bl_int_19_108 bl_int_18_108 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c109
+ bl_int_19_109 bl_int_18_109 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c110
+ bl_int_19_110 bl_int_18_110 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c111
+ bl_int_19_111 bl_int_18_111 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c112
+ bl_int_19_112 bl_int_18_112 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c113
+ bl_int_19_113 bl_int_18_113 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c114
+ bl_int_19_114 bl_int_18_114 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c115
+ bl_int_19_115 bl_int_18_115 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c116
+ bl_int_19_116 bl_int_18_116 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c117
+ bl_int_19_117 bl_int_18_117 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c118
+ bl_int_19_118 bl_int_18_118 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c119
+ bl_int_19_119 bl_int_18_119 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c120
+ bl_int_19_120 bl_int_18_120 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c121
+ bl_int_19_121 bl_int_18_121 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c122
+ bl_int_19_122 bl_int_18_122 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c123
+ bl_int_19_123 bl_int_18_123 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c124
+ bl_int_19_124 bl_int_18_124 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c125
+ bl_int_19_125 bl_int_18_125 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c126
+ bl_int_19_126 bl_int_18_126 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c127
+ bl_int_19_127 bl_int_18_127 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c128
+ bl_int_19_128 bl_int_18_128 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c129
+ bl_int_19_129 bl_int_18_129 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c130
+ bl_int_19_130 bl_int_18_130 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c131
+ bl_int_19_131 bl_int_18_131 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c132
+ bl_int_19_132 bl_int_18_132 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c133
+ bl_int_19_133 bl_int_18_133 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c134
+ bl_int_19_134 bl_int_18_134 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c135
+ bl_int_19_135 bl_int_18_135 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c136
+ bl_int_19_136 bl_int_18_136 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c137
+ bl_int_19_137 bl_int_18_137 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c138
+ bl_int_19_138 bl_int_18_138 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c139
+ bl_int_19_139 bl_int_18_139 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c140
+ bl_int_19_140 bl_int_18_140 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c141
+ bl_int_19_141 bl_int_18_141 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c142
+ bl_int_19_142 bl_int_18_142 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c143
+ bl_int_19_143 bl_int_18_143 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c144
+ bl_int_19_144 bl_int_18_144 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c145
+ bl_int_19_145 bl_int_18_145 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c146
+ bl_int_19_146 bl_int_18_146 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c147
+ bl_int_19_147 bl_int_18_147 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c148
+ bl_int_19_148 bl_int_18_148 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c149
+ bl_int_19_149 bl_int_18_149 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c150
+ bl_int_19_150 bl_int_18_150 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c151
+ bl_int_19_151 bl_int_18_151 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c152
+ bl_int_19_152 bl_int_18_152 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c153
+ bl_int_19_153 bl_int_18_153 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c154
+ bl_int_19_154 bl_int_18_154 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c155
+ bl_int_19_155 bl_int_18_155 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c156
+ bl_int_19_156 bl_int_18_156 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c157
+ bl_int_19_157 bl_int_18_157 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c158
+ bl_int_19_158 bl_int_18_158 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c159
+ bl_int_19_159 bl_int_18_159 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c160
+ bl_int_19_160 bl_int_18_160 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c161
+ bl_int_19_161 bl_int_18_161 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c162
+ bl_int_19_162 bl_int_18_162 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c163
+ bl_int_19_163 bl_int_18_163 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c164
+ bl_int_19_164 bl_int_18_164 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c165
+ bl_int_19_165 bl_int_18_165 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c166
+ bl_int_19_166 bl_int_18_166 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c167
+ bl_int_19_167 bl_int_18_167 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c168
+ bl_int_19_168 bl_int_18_168 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c169
+ bl_int_19_169 bl_int_18_169 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c170
+ bl_int_19_170 bl_int_18_170 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c171
+ bl_int_19_171 bl_int_18_171 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c172
+ bl_int_19_172 bl_int_18_172 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c173
+ bl_int_19_173 bl_int_18_173 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c174
+ bl_int_19_174 bl_int_18_174 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c175
+ bl_int_19_175 bl_int_18_175 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c176
+ bl_int_19_176 bl_int_18_176 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c177
+ bl_int_19_177 bl_int_18_177 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c178
+ bl_int_19_178 bl_int_18_178 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c179
+ bl_int_19_179 bl_int_18_179 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c180
+ bl_int_19_180 bl_int_18_180 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c181
+ bl_int_19_181 bl_int_18_181 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c182
+ bl_int_19_182 bl_int_18_182 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r19_c183
+ bl_int_19_183 bl_int_18_183 wl_0_19 gnd
+ sram_rom_base_one_cell
Xbit_r20_c0
+ bl_int_20_0 bl_int_19_0 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c1
+ bl_int_20_1 bl_int_19_1 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c2
+ bl_int_20_2 bl_int_19_2 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c3
+ bl_int_20_3 bl_int_19_3 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c4
+ bl_int_20_4 bl_int_19_4 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c5
+ bl_int_20_5 bl_int_19_5 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c6
+ bl_int_20_6 bl_int_19_6 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c7
+ bl_int_20_7 bl_int_19_7 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c8
+ bl_int_20_8 bl_int_19_8 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c9
+ bl_int_20_9 bl_int_19_9 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c10
+ bl_int_20_10 bl_int_19_10 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c11
+ bl_int_20_11 bl_int_19_11 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c12
+ bl_int_20_12 bl_int_19_12 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c13
+ bl_int_20_13 bl_int_19_13 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c14
+ bl_int_20_14 bl_int_19_14 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c15
+ bl_int_20_15 bl_int_19_15 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c16
+ bl_int_20_16 bl_int_19_16 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c17
+ bl_int_20_17 bl_int_19_17 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c18
+ bl_int_20_18 bl_int_19_18 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c19
+ bl_int_20_19 bl_int_19_19 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c20
+ bl_int_20_20 bl_int_19_20 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c21
+ bl_int_20_21 bl_int_19_21 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c22
+ bl_int_20_22 bl_int_19_22 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c23
+ bl_int_20_23 bl_int_19_23 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c24
+ bl_int_20_24 bl_int_19_24 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c25
+ bl_int_20_25 bl_int_19_25 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c26
+ bl_int_20_26 bl_int_19_26 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c27
+ bl_int_20_27 bl_int_19_27 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c28
+ bl_int_20_28 bl_int_19_28 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c29
+ bl_int_20_29 bl_int_19_29 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c30
+ bl_int_20_30 bl_int_19_30 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c31
+ bl_int_20_31 bl_int_19_31 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c32
+ bl_int_20_32 bl_int_19_32 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c33
+ bl_int_20_33 bl_int_19_33 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c34
+ bl_int_20_34 bl_int_19_34 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c35
+ bl_int_20_35 bl_int_19_35 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c36
+ bl_int_20_36 bl_int_19_36 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c37
+ bl_int_20_37 bl_int_19_37 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c38
+ bl_int_20_38 bl_int_19_38 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c39
+ bl_int_20_39 bl_int_19_39 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c40
+ bl_int_20_40 bl_int_19_40 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c41
+ bl_int_20_41 bl_int_19_41 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c42
+ bl_int_20_42 bl_int_19_42 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c43
+ bl_int_20_43 bl_int_19_43 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c44
+ bl_int_20_44 bl_int_19_44 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c45
+ bl_int_20_45 bl_int_19_45 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c46
+ bl_int_20_46 bl_int_19_46 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c47
+ bl_int_20_47 bl_int_19_47 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c48
+ bl_int_20_48 bl_int_19_48 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c49
+ bl_int_20_49 bl_int_19_49 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c50
+ bl_int_20_50 bl_int_19_50 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c51
+ bl_int_20_51 bl_int_19_51 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c52
+ bl_int_20_52 bl_int_19_52 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c53
+ bl_int_20_53 bl_int_19_53 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c54
+ bl_int_20_54 bl_int_19_54 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c55
+ bl_int_20_55 bl_int_19_55 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c56
+ bl_int_20_56 bl_int_19_56 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c57
+ bl_int_20_57 bl_int_19_57 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c58
+ bl_int_20_58 bl_int_19_58 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c59
+ bl_int_20_59 bl_int_19_59 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c60
+ bl_int_20_60 bl_int_19_60 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c61
+ bl_int_20_61 bl_int_19_61 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c62
+ bl_int_20_62 bl_int_19_62 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c63
+ bl_int_20_63 bl_int_19_63 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c64
+ bl_int_20_64 bl_int_19_64 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c65
+ bl_int_20_65 bl_int_19_65 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c66
+ bl_int_20_66 bl_int_19_66 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c67
+ bl_int_20_67 bl_int_19_67 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c68
+ bl_int_20_68 bl_int_19_68 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c69
+ bl_int_20_69 bl_int_19_69 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c70
+ bl_int_20_70 bl_int_19_70 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c71
+ bl_int_20_71 bl_int_19_71 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c72
+ bl_int_20_72 bl_int_19_72 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c73
+ bl_int_20_73 bl_int_19_73 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c74
+ bl_int_20_74 bl_int_19_74 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c75
+ bl_int_20_75 bl_int_19_75 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c76
+ bl_int_20_76 bl_int_19_76 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c77
+ bl_int_20_77 bl_int_19_77 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c78
+ bl_int_20_78 bl_int_19_78 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c79
+ bl_int_20_79 bl_int_19_79 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c80
+ bl_int_20_80 bl_int_19_80 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c81
+ bl_int_20_81 bl_int_19_81 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c82
+ bl_int_20_82 bl_int_19_82 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c83
+ bl_int_20_83 bl_int_19_83 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c84
+ bl_int_20_84 bl_int_19_84 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c85
+ bl_int_20_85 bl_int_19_85 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c86
+ bl_int_20_86 bl_int_19_86 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c87
+ bl_int_20_87 bl_int_19_87 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c88
+ bl_int_20_88 bl_int_19_88 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c89
+ bl_int_20_89 bl_int_19_89 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c90
+ bl_int_20_90 bl_int_19_90 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c91
+ bl_int_20_91 bl_int_19_91 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c92
+ bl_int_20_92 bl_int_19_92 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c93
+ bl_int_20_93 bl_int_19_93 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c94
+ bl_int_20_94 bl_int_19_94 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c95
+ bl_int_20_95 bl_int_19_95 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c96
+ bl_int_20_96 bl_int_19_96 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c97
+ bl_int_20_97 bl_int_19_97 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c98
+ bl_int_20_98 bl_int_19_98 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c99
+ bl_int_20_99 bl_int_19_99 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c100
+ bl_int_20_100 bl_int_19_100 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c101
+ bl_int_20_101 bl_int_19_101 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c102
+ bl_int_20_102 bl_int_19_102 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c103
+ bl_int_20_103 bl_int_19_103 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c104
+ bl_int_20_104 bl_int_19_104 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c105
+ bl_int_20_105 bl_int_19_105 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c106
+ bl_int_20_106 bl_int_19_106 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c107
+ bl_int_20_107 bl_int_19_107 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c108
+ bl_int_20_108 bl_int_19_108 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c109
+ bl_int_20_109 bl_int_19_109 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c110
+ bl_int_20_110 bl_int_19_110 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c111
+ bl_int_20_111 bl_int_19_111 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c112
+ bl_int_20_112 bl_int_19_112 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c113
+ bl_int_20_113 bl_int_19_113 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c114
+ bl_int_20_114 bl_int_19_114 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c115
+ bl_int_20_115 bl_int_19_115 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c116
+ bl_int_20_116 bl_int_19_116 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c117
+ bl_int_20_117 bl_int_19_117 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c118
+ bl_int_20_118 bl_int_19_118 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c119
+ bl_int_20_119 bl_int_19_119 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c120
+ bl_int_20_120 bl_int_19_120 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c121
+ bl_int_20_121 bl_int_19_121 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c122
+ bl_int_20_122 bl_int_19_122 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c123
+ bl_int_20_123 bl_int_19_123 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c124
+ bl_int_20_124 bl_int_19_124 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c125
+ bl_int_20_125 bl_int_19_125 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c126
+ bl_int_20_126 bl_int_19_126 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c127
+ bl_int_20_127 bl_int_19_127 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c128
+ bl_int_20_128 bl_int_19_128 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c129
+ bl_int_20_129 bl_int_19_129 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c130
+ bl_int_20_130 bl_int_19_130 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c131
+ bl_int_20_131 bl_int_19_131 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c132
+ bl_int_20_132 bl_int_19_132 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c133
+ bl_int_20_133 bl_int_19_133 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c134
+ bl_int_20_134 bl_int_19_134 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c135
+ bl_int_20_135 bl_int_19_135 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c136
+ bl_int_20_136 bl_int_19_136 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c137
+ bl_int_20_137 bl_int_19_137 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c138
+ bl_int_20_138 bl_int_19_138 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c139
+ bl_int_20_139 bl_int_19_139 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c140
+ bl_int_20_140 bl_int_19_140 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c141
+ bl_int_20_141 bl_int_19_141 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c142
+ bl_int_20_142 bl_int_19_142 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c143
+ bl_int_20_143 bl_int_19_143 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c144
+ bl_int_20_144 bl_int_19_144 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c145
+ bl_int_20_145 bl_int_19_145 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c146
+ bl_int_20_146 bl_int_19_146 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c147
+ bl_int_20_147 bl_int_19_147 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c148
+ bl_int_20_148 bl_int_19_148 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c149
+ bl_int_20_149 bl_int_19_149 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c150
+ bl_int_20_150 bl_int_19_150 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c151
+ bl_int_20_151 bl_int_19_151 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c152
+ bl_int_20_152 bl_int_19_152 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c153
+ bl_int_20_153 bl_int_19_153 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c154
+ bl_int_20_154 bl_int_19_154 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c155
+ bl_int_20_155 bl_int_19_155 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c156
+ bl_int_20_156 bl_int_19_156 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c157
+ bl_int_20_157 bl_int_19_157 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c158
+ bl_int_20_158 bl_int_19_158 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c159
+ bl_int_20_159 bl_int_19_159 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c160
+ bl_int_20_160 bl_int_19_160 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c161
+ bl_int_20_161 bl_int_19_161 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c162
+ bl_int_20_162 bl_int_19_162 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c163
+ bl_int_20_163 bl_int_19_163 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c164
+ bl_int_20_164 bl_int_19_164 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c165
+ bl_int_20_165 bl_int_19_165 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c166
+ bl_int_20_166 bl_int_19_166 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c167
+ bl_int_20_167 bl_int_19_167 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c168
+ bl_int_20_168 bl_int_19_168 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c169
+ bl_int_20_169 bl_int_19_169 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c170
+ bl_int_20_170 bl_int_19_170 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c171
+ bl_int_20_171 bl_int_19_171 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c172
+ bl_int_20_172 bl_int_19_172 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c173
+ bl_int_20_173 bl_int_19_173 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c174
+ bl_int_20_174 bl_int_19_174 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c175
+ bl_int_20_175 bl_int_19_175 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c176
+ bl_int_20_176 bl_int_19_176 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c177
+ bl_int_20_177 bl_int_19_177 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c178
+ bl_int_20_178 bl_int_19_178 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c179
+ bl_int_20_179 bl_int_19_179 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c180
+ bl_int_20_180 bl_int_19_180 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c181
+ bl_int_20_181 bl_int_19_181 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c182
+ bl_int_20_182 bl_int_19_182 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r20_c183
+ bl_int_20_183 bl_int_19_183 wl_0_20 gnd
+ sram_rom_base_one_cell
Xbit_r21_c0
+ bl_int_21_0 bl_int_20_0 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c1
+ bl_int_21_1 bl_int_20_1 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c2
+ bl_int_21_2 bl_int_20_2 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c3
+ bl_int_21_3 bl_int_20_3 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c4
+ bl_int_21_4 bl_int_20_4 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c5
+ bl_int_21_5 bl_int_20_5 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c6
+ bl_int_21_6 bl_int_20_6 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c7
+ bl_int_21_7 bl_int_20_7 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c8
+ bl_int_21_8 bl_int_20_8 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c9
+ bl_int_21_9 bl_int_20_9 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c10
+ bl_int_21_10 bl_int_20_10 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c11
+ bl_int_21_11 bl_int_20_11 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c12
+ bl_int_21_12 bl_int_20_12 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c13
+ bl_int_21_13 bl_int_20_13 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c14
+ bl_int_21_14 bl_int_20_14 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c15
+ bl_int_21_15 bl_int_20_15 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c16
+ bl_int_21_16 bl_int_20_16 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c17
+ bl_int_21_17 bl_int_20_17 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c18
+ bl_int_21_18 bl_int_20_18 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c19
+ bl_int_21_19 bl_int_20_19 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c20
+ bl_int_21_20 bl_int_20_20 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c21
+ bl_int_21_21 bl_int_20_21 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c22
+ bl_int_21_22 bl_int_20_22 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c23
+ bl_int_21_23 bl_int_20_23 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c24
+ bl_int_21_24 bl_int_20_24 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c25
+ bl_int_21_25 bl_int_20_25 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c26
+ bl_int_21_26 bl_int_20_26 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c27
+ bl_int_21_27 bl_int_20_27 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c28
+ bl_int_21_28 bl_int_20_28 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c29
+ bl_int_21_29 bl_int_20_29 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c30
+ bl_int_21_30 bl_int_20_30 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c31
+ bl_int_21_31 bl_int_20_31 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c32
+ bl_int_21_32 bl_int_20_32 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c33
+ bl_int_21_33 bl_int_20_33 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c34
+ bl_int_21_34 bl_int_20_34 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c35
+ bl_int_21_35 bl_int_20_35 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c36
+ bl_int_21_36 bl_int_20_36 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c37
+ bl_int_21_37 bl_int_20_37 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c38
+ bl_int_21_38 bl_int_20_38 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c39
+ bl_int_21_39 bl_int_20_39 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c40
+ bl_int_21_40 bl_int_20_40 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c41
+ bl_int_21_41 bl_int_20_41 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c42
+ bl_int_21_42 bl_int_20_42 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c43
+ bl_int_21_43 bl_int_20_43 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c44
+ bl_int_21_44 bl_int_20_44 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c45
+ bl_int_21_45 bl_int_20_45 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c46
+ bl_int_21_46 bl_int_20_46 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c47
+ bl_int_21_47 bl_int_20_47 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c48
+ bl_int_21_48 bl_int_20_48 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c49
+ bl_int_21_49 bl_int_20_49 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c50
+ bl_int_21_50 bl_int_20_50 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c51
+ bl_int_21_51 bl_int_20_51 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c52
+ bl_int_21_52 bl_int_20_52 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c53
+ bl_int_21_53 bl_int_20_53 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c54
+ bl_int_21_54 bl_int_20_54 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c55
+ bl_int_21_55 bl_int_20_55 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c56
+ bl_int_21_56 bl_int_20_56 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c57
+ bl_int_21_57 bl_int_20_57 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c58
+ bl_int_21_58 bl_int_20_58 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c59
+ bl_int_21_59 bl_int_20_59 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c60
+ bl_int_21_60 bl_int_20_60 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c61
+ bl_int_21_61 bl_int_20_61 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c62
+ bl_int_21_62 bl_int_20_62 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c63
+ bl_int_21_63 bl_int_20_63 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c64
+ bl_int_21_64 bl_int_20_64 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c65
+ bl_int_21_65 bl_int_20_65 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c66
+ bl_int_21_66 bl_int_20_66 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c67
+ bl_int_21_67 bl_int_20_67 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c68
+ bl_int_21_68 bl_int_20_68 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c69
+ bl_int_21_69 bl_int_20_69 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c70
+ bl_int_21_70 bl_int_20_70 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c71
+ bl_int_21_71 bl_int_20_71 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c72
+ bl_int_21_72 bl_int_20_72 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c73
+ bl_int_21_73 bl_int_20_73 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c74
+ bl_int_21_74 bl_int_20_74 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c75
+ bl_int_21_75 bl_int_20_75 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c76
+ bl_int_21_76 bl_int_20_76 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c77
+ bl_int_21_77 bl_int_20_77 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c78
+ bl_int_21_78 bl_int_20_78 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c79
+ bl_int_21_79 bl_int_20_79 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c80
+ bl_int_21_80 bl_int_20_80 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c81
+ bl_int_21_81 bl_int_20_81 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c82
+ bl_int_21_82 bl_int_20_82 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c83
+ bl_int_21_83 bl_int_20_83 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c84
+ bl_int_21_84 bl_int_20_84 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c85
+ bl_int_21_85 bl_int_20_85 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c86
+ bl_int_21_86 bl_int_20_86 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c87
+ bl_int_21_87 bl_int_20_87 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c88
+ bl_int_21_88 bl_int_20_88 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c89
+ bl_int_21_89 bl_int_20_89 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c90
+ bl_int_21_90 bl_int_20_90 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c91
+ bl_int_21_91 bl_int_20_91 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c92
+ bl_int_21_92 bl_int_20_92 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c93
+ bl_int_21_93 bl_int_20_93 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c94
+ bl_int_21_94 bl_int_20_94 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c95
+ bl_int_21_95 bl_int_20_95 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c96
+ bl_int_21_96 bl_int_20_96 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c97
+ bl_int_21_97 bl_int_20_97 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c98
+ bl_int_21_98 bl_int_20_98 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c99
+ bl_int_21_99 bl_int_20_99 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c100
+ bl_int_21_100 bl_int_20_100 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c101
+ bl_int_21_101 bl_int_20_101 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c102
+ bl_int_21_102 bl_int_20_102 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c103
+ bl_int_21_103 bl_int_20_103 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c104
+ bl_int_21_104 bl_int_20_104 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c105
+ bl_int_21_105 bl_int_20_105 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c106
+ bl_int_21_106 bl_int_20_106 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c107
+ bl_int_21_107 bl_int_20_107 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c108
+ bl_int_21_108 bl_int_20_108 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c109
+ bl_int_21_109 bl_int_20_109 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c110
+ bl_int_21_110 bl_int_20_110 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c111
+ bl_int_21_111 bl_int_20_111 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c112
+ bl_int_21_112 bl_int_20_112 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c113
+ bl_int_21_113 bl_int_20_113 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c114
+ bl_int_21_114 bl_int_20_114 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c115
+ bl_int_21_115 bl_int_20_115 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c116
+ bl_int_21_116 bl_int_20_116 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c117
+ bl_int_21_117 bl_int_20_117 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c118
+ bl_int_21_118 bl_int_20_118 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c119
+ bl_int_21_119 bl_int_20_119 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c120
+ bl_int_21_120 bl_int_20_120 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c121
+ bl_int_21_121 bl_int_20_121 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c122
+ bl_int_21_122 bl_int_20_122 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c123
+ bl_int_21_123 bl_int_20_123 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c124
+ bl_int_21_124 bl_int_20_124 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c125
+ bl_int_21_125 bl_int_20_125 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c126
+ bl_int_21_126 bl_int_20_126 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c127
+ bl_int_21_127 bl_int_20_127 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c128
+ bl_int_21_128 bl_int_20_128 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c129
+ bl_int_21_129 bl_int_20_129 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c130
+ bl_int_21_130 bl_int_20_130 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c131
+ bl_int_21_131 bl_int_20_131 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c132
+ bl_int_21_132 bl_int_20_132 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c133
+ bl_int_21_133 bl_int_20_133 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c134
+ bl_int_21_134 bl_int_20_134 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c135
+ bl_int_21_135 bl_int_20_135 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c136
+ bl_int_21_136 bl_int_20_136 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c137
+ bl_int_21_137 bl_int_20_137 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c138
+ bl_int_21_138 bl_int_20_138 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c139
+ bl_int_21_139 bl_int_20_139 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c140
+ bl_int_21_140 bl_int_20_140 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c141
+ bl_int_21_141 bl_int_20_141 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c142
+ bl_int_21_142 bl_int_20_142 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c143
+ bl_int_21_143 bl_int_20_143 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c144
+ bl_int_21_144 bl_int_20_144 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c145
+ bl_int_21_145 bl_int_20_145 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c146
+ bl_int_21_146 bl_int_20_146 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c147
+ bl_int_21_147 bl_int_20_147 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c148
+ bl_int_21_148 bl_int_20_148 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c149
+ bl_int_21_149 bl_int_20_149 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c150
+ bl_int_21_150 bl_int_20_150 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c151
+ bl_int_21_151 bl_int_20_151 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c152
+ bl_int_21_152 bl_int_20_152 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c153
+ bl_int_21_153 bl_int_20_153 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c154
+ bl_int_21_154 bl_int_20_154 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c155
+ bl_int_21_155 bl_int_20_155 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c156
+ bl_int_21_156 bl_int_20_156 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c157
+ bl_int_21_157 bl_int_20_157 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c158
+ bl_int_21_158 bl_int_20_158 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c159
+ bl_int_21_159 bl_int_20_159 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c160
+ bl_int_21_160 bl_int_20_160 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c161
+ bl_int_21_161 bl_int_20_161 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c162
+ bl_int_21_162 bl_int_20_162 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c163
+ bl_int_21_163 bl_int_20_163 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c164
+ bl_int_21_164 bl_int_20_164 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c165
+ bl_int_21_165 bl_int_20_165 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c166
+ bl_int_21_166 bl_int_20_166 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c167
+ bl_int_21_167 bl_int_20_167 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c168
+ bl_int_21_168 bl_int_20_168 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c169
+ bl_int_21_169 bl_int_20_169 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c170
+ bl_int_21_170 bl_int_20_170 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c171
+ bl_int_21_171 bl_int_20_171 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c172
+ bl_int_21_172 bl_int_20_172 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c173
+ bl_int_21_173 bl_int_20_173 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c174
+ bl_int_21_174 bl_int_20_174 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c175
+ bl_int_21_175 bl_int_20_175 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c176
+ bl_int_21_176 bl_int_20_176 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c177
+ bl_int_21_177 bl_int_20_177 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c178
+ bl_int_21_178 bl_int_20_178 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c179
+ bl_int_21_179 bl_int_20_179 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c180
+ bl_int_21_180 bl_int_20_180 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c181
+ bl_int_21_181 bl_int_20_181 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c182
+ bl_int_21_182 bl_int_20_182 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r21_c183
+ bl_int_21_183 bl_int_20_183 wl_0_21 gnd
+ sram_rom_base_one_cell
Xbit_r22_c0
+ bl_int_22_0 bl_int_21_0 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c1
+ bl_int_22_1 bl_int_21_1 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c2
+ bl_int_22_2 bl_int_21_2 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c3
+ bl_int_22_3 bl_int_21_3 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c4
+ bl_int_22_4 bl_int_21_4 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c5
+ bl_int_22_5 bl_int_21_5 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c6
+ bl_int_22_6 bl_int_21_6 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c7
+ bl_int_22_7 bl_int_21_7 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c8
+ bl_int_22_8 bl_int_21_8 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c9
+ bl_int_22_9 bl_int_21_9 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c10
+ bl_int_22_10 bl_int_21_10 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c11
+ bl_int_22_11 bl_int_21_11 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c12
+ bl_int_22_12 bl_int_21_12 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c13
+ bl_int_22_13 bl_int_21_13 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c14
+ bl_int_22_14 bl_int_21_14 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c15
+ bl_int_22_15 bl_int_21_15 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c16
+ bl_int_22_16 bl_int_21_16 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c17
+ bl_int_22_17 bl_int_21_17 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c18
+ bl_int_22_18 bl_int_21_18 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c19
+ bl_int_22_19 bl_int_21_19 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c20
+ bl_int_22_20 bl_int_21_20 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c21
+ bl_int_22_21 bl_int_21_21 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c22
+ bl_int_22_22 bl_int_21_22 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c23
+ bl_int_22_23 bl_int_21_23 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c24
+ bl_int_22_24 bl_int_21_24 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c25
+ bl_int_22_25 bl_int_21_25 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c26
+ bl_int_22_26 bl_int_21_26 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c27
+ bl_int_22_27 bl_int_21_27 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c28
+ bl_int_22_28 bl_int_21_28 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c29
+ bl_int_22_29 bl_int_21_29 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c30
+ bl_int_22_30 bl_int_21_30 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c31
+ bl_int_22_31 bl_int_21_31 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c32
+ bl_int_22_32 bl_int_21_32 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c33
+ bl_int_22_33 bl_int_21_33 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c34
+ bl_int_22_34 bl_int_21_34 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c35
+ bl_int_22_35 bl_int_21_35 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c36
+ bl_int_22_36 bl_int_21_36 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c37
+ bl_int_22_37 bl_int_21_37 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c38
+ bl_int_22_38 bl_int_21_38 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c39
+ bl_int_22_39 bl_int_21_39 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c40
+ bl_int_22_40 bl_int_21_40 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c41
+ bl_int_22_41 bl_int_21_41 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c42
+ bl_int_22_42 bl_int_21_42 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c43
+ bl_int_22_43 bl_int_21_43 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c44
+ bl_int_22_44 bl_int_21_44 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c45
+ bl_int_22_45 bl_int_21_45 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c46
+ bl_int_22_46 bl_int_21_46 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c47
+ bl_int_22_47 bl_int_21_47 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c48
+ bl_int_22_48 bl_int_21_48 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c49
+ bl_int_22_49 bl_int_21_49 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c50
+ bl_int_22_50 bl_int_21_50 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c51
+ bl_int_22_51 bl_int_21_51 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c52
+ bl_int_22_52 bl_int_21_52 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c53
+ bl_int_22_53 bl_int_21_53 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c54
+ bl_int_22_54 bl_int_21_54 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c55
+ bl_int_22_55 bl_int_21_55 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c56
+ bl_int_22_56 bl_int_21_56 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c57
+ bl_int_22_57 bl_int_21_57 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c58
+ bl_int_22_58 bl_int_21_58 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c59
+ bl_int_22_59 bl_int_21_59 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c60
+ bl_int_22_60 bl_int_21_60 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c61
+ bl_int_22_61 bl_int_21_61 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c62
+ bl_int_22_62 bl_int_21_62 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c63
+ bl_int_22_63 bl_int_21_63 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c64
+ bl_int_22_64 bl_int_21_64 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c65
+ bl_int_22_65 bl_int_21_65 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c66
+ bl_int_22_66 bl_int_21_66 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c67
+ bl_int_22_67 bl_int_21_67 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c68
+ bl_int_22_68 bl_int_21_68 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c69
+ bl_int_22_69 bl_int_21_69 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c70
+ bl_int_22_70 bl_int_21_70 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c71
+ bl_int_22_71 bl_int_21_71 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c72
+ bl_int_22_72 bl_int_21_72 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c73
+ bl_int_22_73 bl_int_21_73 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c74
+ bl_int_22_74 bl_int_21_74 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c75
+ bl_int_22_75 bl_int_21_75 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c76
+ bl_int_22_76 bl_int_21_76 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c77
+ bl_int_22_77 bl_int_21_77 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c78
+ bl_int_22_78 bl_int_21_78 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c79
+ bl_int_22_79 bl_int_21_79 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c80
+ bl_int_22_80 bl_int_21_80 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c81
+ bl_int_22_81 bl_int_21_81 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c82
+ bl_int_22_82 bl_int_21_82 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c83
+ bl_int_22_83 bl_int_21_83 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c84
+ bl_int_22_84 bl_int_21_84 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c85
+ bl_int_22_85 bl_int_21_85 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c86
+ bl_int_22_86 bl_int_21_86 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c87
+ bl_int_22_87 bl_int_21_87 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c88
+ bl_int_22_88 bl_int_21_88 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c89
+ bl_int_22_89 bl_int_21_89 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c90
+ bl_int_22_90 bl_int_21_90 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c91
+ bl_int_22_91 bl_int_21_91 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c92
+ bl_int_22_92 bl_int_21_92 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c93
+ bl_int_22_93 bl_int_21_93 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c94
+ bl_int_22_94 bl_int_21_94 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c95
+ bl_int_22_95 bl_int_21_95 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c96
+ bl_int_22_96 bl_int_21_96 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c97
+ bl_int_22_97 bl_int_21_97 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c98
+ bl_int_22_98 bl_int_21_98 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c99
+ bl_int_22_99 bl_int_21_99 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c100
+ bl_int_22_100 bl_int_21_100 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c101
+ bl_int_22_101 bl_int_21_101 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c102
+ bl_int_22_102 bl_int_21_102 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c103
+ bl_int_22_103 bl_int_21_103 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c104
+ bl_int_22_104 bl_int_21_104 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c105
+ bl_int_22_105 bl_int_21_105 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c106
+ bl_int_22_106 bl_int_21_106 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c107
+ bl_int_22_107 bl_int_21_107 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c108
+ bl_int_22_108 bl_int_21_108 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c109
+ bl_int_22_109 bl_int_21_109 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c110
+ bl_int_22_110 bl_int_21_110 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c111
+ bl_int_22_111 bl_int_21_111 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c112
+ bl_int_22_112 bl_int_21_112 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c113
+ bl_int_22_113 bl_int_21_113 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c114
+ bl_int_22_114 bl_int_21_114 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c115
+ bl_int_22_115 bl_int_21_115 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c116
+ bl_int_22_116 bl_int_21_116 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c117
+ bl_int_22_117 bl_int_21_117 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c118
+ bl_int_22_118 bl_int_21_118 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c119
+ bl_int_22_119 bl_int_21_119 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c120
+ bl_int_22_120 bl_int_21_120 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c121
+ bl_int_22_121 bl_int_21_121 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c122
+ bl_int_22_122 bl_int_21_122 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c123
+ bl_int_22_123 bl_int_21_123 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c124
+ bl_int_22_124 bl_int_21_124 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c125
+ bl_int_22_125 bl_int_21_125 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c126
+ bl_int_22_126 bl_int_21_126 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c127
+ bl_int_22_127 bl_int_21_127 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c128
+ bl_int_22_128 bl_int_21_128 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c129
+ bl_int_22_129 bl_int_21_129 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c130
+ bl_int_22_130 bl_int_21_130 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c131
+ bl_int_22_131 bl_int_21_131 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c132
+ bl_int_22_132 bl_int_21_132 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c133
+ bl_int_22_133 bl_int_21_133 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c134
+ bl_int_22_134 bl_int_21_134 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c135
+ bl_int_22_135 bl_int_21_135 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c136
+ bl_int_22_136 bl_int_21_136 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c137
+ bl_int_22_137 bl_int_21_137 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c138
+ bl_int_22_138 bl_int_21_138 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c139
+ bl_int_22_139 bl_int_21_139 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c140
+ bl_int_22_140 bl_int_21_140 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c141
+ bl_int_22_141 bl_int_21_141 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c142
+ bl_int_22_142 bl_int_21_142 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c143
+ bl_int_22_143 bl_int_21_143 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c144
+ bl_int_22_144 bl_int_21_144 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c145
+ bl_int_22_145 bl_int_21_145 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c146
+ bl_int_22_146 bl_int_21_146 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c147
+ bl_int_22_147 bl_int_21_147 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c148
+ bl_int_22_148 bl_int_21_148 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c149
+ bl_int_22_149 bl_int_21_149 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c150
+ bl_int_22_150 bl_int_21_150 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c151
+ bl_int_22_151 bl_int_21_151 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c152
+ bl_int_22_152 bl_int_21_152 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c153
+ bl_int_22_153 bl_int_21_153 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c154
+ bl_int_22_154 bl_int_21_154 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c155
+ bl_int_22_155 bl_int_21_155 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c156
+ bl_int_22_156 bl_int_21_156 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c157
+ bl_int_22_157 bl_int_21_157 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c158
+ bl_int_22_158 bl_int_21_158 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c159
+ bl_int_22_159 bl_int_21_159 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c160
+ bl_int_22_160 bl_int_21_160 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c161
+ bl_int_22_161 bl_int_21_161 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c162
+ bl_int_22_162 bl_int_21_162 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c163
+ bl_int_22_163 bl_int_21_163 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c164
+ bl_int_22_164 bl_int_21_164 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c165
+ bl_int_22_165 bl_int_21_165 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c166
+ bl_int_22_166 bl_int_21_166 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c167
+ bl_int_22_167 bl_int_21_167 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c168
+ bl_int_22_168 bl_int_21_168 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c169
+ bl_int_22_169 bl_int_21_169 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c170
+ bl_int_22_170 bl_int_21_170 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c171
+ bl_int_22_171 bl_int_21_171 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c172
+ bl_int_22_172 bl_int_21_172 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c173
+ bl_int_22_173 bl_int_21_173 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c174
+ bl_int_22_174 bl_int_21_174 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c175
+ bl_int_22_175 bl_int_21_175 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c176
+ bl_int_22_176 bl_int_21_176 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c177
+ bl_int_22_177 bl_int_21_177 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c178
+ bl_int_22_178 bl_int_21_178 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c179
+ bl_int_22_179 bl_int_21_179 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c180
+ bl_int_22_180 bl_int_21_180 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c181
+ bl_int_22_181 bl_int_21_181 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c182
+ bl_int_22_182 bl_int_21_182 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r22_c183
+ bl_int_22_183 bl_int_21_183 wl_0_22 gnd
+ sram_rom_base_one_cell
Xbit_r23_c0
+ bl_int_23_0 bl_int_22_0 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c1
+ bl_int_23_1 bl_int_22_1 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c2
+ bl_int_23_2 bl_int_22_2 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c3
+ bl_int_23_3 bl_int_22_3 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c4
+ bl_int_23_4 bl_int_22_4 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c5
+ bl_int_23_5 bl_int_22_5 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c6
+ bl_int_23_6 bl_int_22_6 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c7
+ bl_int_23_7 bl_int_22_7 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c8
+ bl_int_23_8 bl_int_22_8 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c9
+ bl_int_23_9 bl_int_22_9 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c10
+ bl_int_23_10 bl_int_22_10 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c11
+ bl_int_23_11 bl_int_22_11 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c12
+ bl_int_23_12 bl_int_22_12 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c13
+ bl_int_23_13 bl_int_22_13 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c14
+ bl_int_23_14 bl_int_22_14 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c15
+ bl_int_23_15 bl_int_22_15 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c16
+ bl_int_23_16 bl_int_22_16 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c17
+ bl_int_23_17 bl_int_22_17 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c18
+ bl_int_23_18 bl_int_22_18 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c19
+ bl_int_23_19 bl_int_22_19 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c20
+ bl_int_23_20 bl_int_22_20 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c21
+ bl_int_23_21 bl_int_22_21 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c22
+ bl_int_23_22 bl_int_22_22 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c23
+ bl_int_23_23 bl_int_22_23 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c24
+ bl_int_23_24 bl_int_22_24 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c25
+ bl_int_23_25 bl_int_22_25 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c26
+ bl_int_23_26 bl_int_22_26 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c27
+ bl_int_23_27 bl_int_22_27 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c28
+ bl_int_23_28 bl_int_22_28 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c29
+ bl_int_23_29 bl_int_22_29 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c30
+ bl_int_23_30 bl_int_22_30 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c31
+ bl_int_23_31 bl_int_22_31 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c32
+ bl_int_23_32 bl_int_22_32 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c33
+ bl_int_23_33 bl_int_22_33 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c34
+ bl_int_23_34 bl_int_22_34 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c35
+ bl_int_23_35 bl_int_22_35 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c36
+ bl_int_23_36 bl_int_22_36 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c37
+ bl_int_23_37 bl_int_22_37 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c38
+ bl_int_23_38 bl_int_22_38 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c39
+ bl_int_23_39 bl_int_22_39 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c40
+ bl_int_23_40 bl_int_22_40 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c41
+ bl_int_23_41 bl_int_22_41 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c42
+ bl_int_23_42 bl_int_22_42 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c43
+ bl_int_23_43 bl_int_22_43 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c44
+ bl_int_23_44 bl_int_22_44 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c45
+ bl_int_23_45 bl_int_22_45 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c46
+ bl_int_23_46 bl_int_22_46 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c47
+ bl_int_23_47 bl_int_22_47 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c48
+ bl_int_23_48 bl_int_22_48 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c49
+ bl_int_23_49 bl_int_22_49 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c50
+ bl_int_23_50 bl_int_22_50 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c51
+ bl_int_23_51 bl_int_22_51 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c52
+ bl_int_23_52 bl_int_22_52 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c53
+ bl_int_23_53 bl_int_22_53 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c54
+ bl_int_23_54 bl_int_22_54 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c55
+ bl_int_23_55 bl_int_22_55 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c56
+ bl_int_23_56 bl_int_22_56 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c57
+ bl_int_23_57 bl_int_22_57 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c58
+ bl_int_23_58 bl_int_22_58 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c59
+ bl_int_23_59 bl_int_22_59 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c60
+ bl_int_23_60 bl_int_22_60 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c61
+ bl_int_23_61 bl_int_22_61 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c62
+ bl_int_23_62 bl_int_22_62 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c63
+ bl_int_23_63 bl_int_22_63 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c64
+ bl_int_23_64 bl_int_22_64 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c65
+ bl_int_23_65 bl_int_22_65 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c66
+ bl_int_23_66 bl_int_22_66 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c67
+ bl_int_23_67 bl_int_22_67 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c68
+ bl_int_23_68 bl_int_22_68 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c69
+ bl_int_23_69 bl_int_22_69 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c70
+ bl_int_23_70 bl_int_22_70 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c71
+ bl_int_23_71 bl_int_22_71 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c72
+ bl_int_23_72 bl_int_22_72 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c73
+ bl_int_23_73 bl_int_22_73 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c74
+ bl_int_23_74 bl_int_22_74 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c75
+ bl_int_23_75 bl_int_22_75 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c76
+ bl_int_23_76 bl_int_22_76 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c77
+ bl_int_23_77 bl_int_22_77 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c78
+ bl_int_23_78 bl_int_22_78 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c79
+ bl_int_23_79 bl_int_22_79 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c80
+ bl_int_23_80 bl_int_22_80 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c81
+ bl_int_23_81 bl_int_22_81 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c82
+ bl_int_23_82 bl_int_22_82 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c83
+ bl_int_23_83 bl_int_22_83 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c84
+ bl_int_23_84 bl_int_22_84 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c85
+ bl_int_23_85 bl_int_22_85 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c86
+ bl_int_23_86 bl_int_22_86 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c87
+ bl_int_23_87 bl_int_22_87 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c88
+ bl_int_23_88 bl_int_22_88 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c89
+ bl_int_23_89 bl_int_22_89 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c90
+ bl_int_23_90 bl_int_22_90 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c91
+ bl_int_23_91 bl_int_22_91 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c92
+ bl_int_23_92 bl_int_22_92 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c93
+ bl_int_23_93 bl_int_22_93 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c94
+ bl_int_23_94 bl_int_22_94 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c95
+ bl_int_23_95 bl_int_22_95 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c96
+ bl_int_23_96 bl_int_22_96 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c97
+ bl_int_23_97 bl_int_22_97 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c98
+ bl_int_23_98 bl_int_22_98 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c99
+ bl_int_23_99 bl_int_22_99 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c100
+ bl_int_23_100 bl_int_22_100 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c101
+ bl_int_23_101 bl_int_22_101 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c102
+ bl_int_23_102 bl_int_22_102 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c103
+ bl_int_23_103 bl_int_22_103 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c104
+ bl_int_23_104 bl_int_22_104 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c105
+ bl_int_23_105 bl_int_22_105 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c106
+ bl_int_23_106 bl_int_22_106 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c107
+ bl_int_23_107 bl_int_22_107 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c108
+ bl_int_23_108 bl_int_22_108 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c109
+ bl_int_23_109 bl_int_22_109 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c110
+ bl_int_23_110 bl_int_22_110 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c111
+ bl_int_23_111 bl_int_22_111 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c112
+ bl_int_23_112 bl_int_22_112 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c113
+ bl_int_23_113 bl_int_22_113 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c114
+ bl_int_23_114 bl_int_22_114 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c115
+ bl_int_23_115 bl_int_22_115 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c116
+ bl_int_23_116 bl_int_22_116 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c117
+ bl_int_23_117 bl_int_22_117 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c118
+ bl_int_23_118 bl_int_22_118 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c119
+ bl_int_23_119 bl_int_22_119 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c120
+ bl_int_23_120 bl_int_22_120 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c121
+ bl_int_23_121 bl_int_22_121 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c122
+ bl_int_23_122 bl_int_22_122 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c123
+ bl_int_23_123 bl_int_22_123 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c124
+ bl_int_23_124 bl_int_22_124 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c125
+ bl_int_23_125 bl_int_22_125 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c126
+ bl_int_23_126 bl_int_22_126 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c127
+ bl_int_23_127 bl_int_22_127 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c128
+ bl_int_23_128 bl_int_22_128 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c129
+ bl_int_23_129 bl_int_22_129 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c130
+ bl_int_23_130 bl_int_22_130 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c131
+ bl_int_23_131 bl_int_22_131 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c132
+ bl_int_23_132 bl_int_22_132 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c133
+ bl_int_23_133 bl_int_22_133 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c134
+ bl_int_23_134 bl_int_22_134 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c135
+ bl_int_23_135 bl_int_22_135 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c136
+ bl_int_23_136 bl_int_22_136 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c137
+ bl_int_23_137 bl_int_22_137 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c138
+ bl_int_23_138 bl_int_22_138 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c139
+ bl_int_23_139 bl_int_22_139 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c140
+ bl_int_23_140 bl_int_22_140 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c141
+ bl_int_23_141 bl_int_22_141 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c142
+ bl_int_23_142 bl_int_22_142 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c143
+ bl_int_23_143 bl_int_22_143 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c144
+ bl_int_23_144 bl_int_22_144 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c145
+ bl_int_23_145 bl_int_22_145 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c146
+ bl_int_23_146 bl_int_22_146 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c147
+ bl_int_23_147 bl_int_22_147 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c148
+ bl_int_23_148 bl_int_22_148 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c149
+ bl_int_23_149 bl_int_22_149 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c150
+ bl_int_23_150 bl_int_22_150 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c151
+ bl_int_23_151 bl_int_22_151 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c152
+ bl_int_23_152 bl_int_22_152 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c153
+ bl_int_23_153 bl_int_22_153 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c154
+ bl_int_23_154 bl_int_22_154 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c155
+ bl_int_23_155 bl_int_22_155 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c156
+ bl_int_23_156 bl_int_22_156 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c157
+ bl_int_23_157 bl_int_22_157 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c158
+ bl_int_23_158 bl_int_22_158 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c159
+ bl_int_23_159 bl_int_22_159 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c160
+ bl_int_23_160 bl_int_22_160 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c161
+ bl_int_23_161 bl_int_22_161 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c162
+ bl_int_23_162 bl_int_22_162 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c163
+ bl_int_23_163 bl_int_22_163 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c164
+ bl_int_23_164 bl_int_22_164 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c165
+ bl_int_23_165 bl_int_22_165 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c166
+ bl_int_23_166 bl_int_22_166 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c167
+ bl_int_23_167 bl_int_22_167 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c168
+ bl_int_23_168 bl_int_22_168 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c169
+ bl_int_23_169 bl_int_22_169 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c170
+ bl_int_23_170 bl_int_22_170 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c171
+ bl_int_23_171 bl_int_22_171 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c172
+ bl_int_23_172 bl_int_22_172 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c173
+ bl_int_23_173 bl_int_22_173 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c174
+ bl_int_23_174 bl_int_22_174 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c175
+ bl_int_23_175 bl_int_22_175 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c176
+ bl_int_23_176 bl_int_22_176 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c177
+ bl_int_23_177 bl_int_22_177 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c178
+ bl_int_23_178 bl_int_22_178 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c179
+ bl_int_23_179 bl_int_22_179 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c180
+ bl_int_23_180 bl_int_22_180 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c181
+ bl_int_23_181 bl_int_22_181 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c182
+ bl_int_23_182 bl_int_22_182 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r23_c183
+ bl_int_23_183 bl_int_22_183 wl_0_23 gnd
+ sram_rom_base_one_cell
Xbit_r24_c0
+ bl_int_24_0 bl_int_23_0 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c1
+ bl_int_24_1 bl_int_23_1 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c2
+ bl_int_24_2 bl_int_23_2 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c3
+ bl_int_24_3 bl_int_23_3 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c4
+ bl_int_24_4 bl_int_23_4 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c5
+ bl_int_24_5 bl_int_23_5 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c6
+ bl_int_24_6 bl_int_23_6 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c7
+ bl_int_24_7 bl_int_23_7 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c8
+ bl_int_24_8 bl_int_23_8 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c9
+ bl_int_24_9 bl_int_23_9 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c10
+ bl_int_24_10 bl_int_23_10 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c11
+ bl_int_24_11 bl_int_23_11 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c12
+ bl_int_24_12 bl_int_23_12 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c13
+ bl_int_24_13 bl_int_23_13 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c14
+ bl_int_24_14 bl_int_23_14 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c15
+ bl_int_24_15 bl_int_23_15 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c16
+ bl_int_24_16 bl_int_23_16 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c17
+ bl_int_24_17 bl_int_23_17 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c18
+ bl_int_24_18 bl_int_23_18 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c19
+ bl_int_24_19 bl_int_23_19 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c20
+ bl_int_24_20 bl_int_23_20 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c21
+ bl_int_24_21 bl_int_23_21 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c22
+ bl_int_24_22 bl_int_23_22 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c23
+ bl_int_24_23 bl_int_23_23 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c24
+ bl_int_24_24 bl_int_23_24 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c25
+ bl_int_24_25 bl_int_23_25 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c26
+ bl_int_24_26 bl_int_23_26 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c27
+ bl_int_24_27 bl_int_23_27 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c28
+ bl_int_24_28 bl_int_23_28 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c29
+ bl_int_24_29 bl_int_23_29 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c30
+ bl_int_24_30 bl_int_23_30 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c31
+ bl_int_24_31 bl_int_23_31 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c32
+ bl_int_24_32 bl_int_23_32 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c33
+ bl_int_24_33 bl_int_23_33 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c34
+ bl_int_24_34 bl_int_23_34 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c35
+ bl_int_24_35 bl_int_23_35 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c36
+ bl_int_24_36 bl_int_23_36 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c37
+ bl_int_24_37 bl_int_23_37 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c38
+ bl_int_24_38 bl_int_23_38 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c39
+ bl_int_24_39 bl_int_23_39 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c40
+ bl_int_24_40 bl_int_23_40 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c41
+ bl_int_24_41 bl_int_23_41 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c42
+ bl_int_24_42 bl_int_23_42 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c43
+ bl_int_24_43 bl_int_23_43 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c44
+ bl_int_24_44 bl_int_23_44 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c45
+ bl_int_24_45 bl_int_23_45 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c46
+ bl_int_24_46 bl_int_23_46 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c47
+ bl_int_24_47 bl_int_23_47 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c48
+ bl_int_24_48 bl_int_23_48 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c49
+ bl_int_24_49 bl_int_23_49 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c50
+ bl_int_24_50 bl_int_23_50 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c51
+ bl_int_24_51 bl_int_23_51 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c52
+ bl_int_24_52 bl_int_23_52 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c53
+ bl_int_24_53 bl_int_23_53 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c54
+ bl_int_24_54 bl_int_23_54 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c55
+ bl_int_24_55 bl_int_23_55 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c56
+ bl_int_24_56 bl_int_23_56 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c57
+ bl_int_24_57 bl_int_23_57 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c58
+ bl_int_24_58 bl_int_23_58 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c59
+ bl_int_24_59 bl_int_23_59 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c60
+ bl_int_24_60 bl_int_23_60 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c61
+ bl_int_24_61 bl_int_23_61 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c62
+ bl_int_24_62 bl_int_23_62 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c63
+ bl_int_24_63 bl_int_23_63 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c64
+ bl_int_24_64 bl_int_23_64 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c65
+ bl_int_24_65 bl_int_23_65 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c66
+ bl_int_24_66 bl_int_23_66 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c67
+ bl_int_24_67 bl_int_23_67 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c68
+ bl_int_24_68 bl_int_23_68 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c69
+ bl_int_24_69 bl_int_23_69 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c70
+ bl_int_24_70 bl_int_23_70 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c71
+ bl_int_24_71 bl_int_23_71 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c72
+ bl_int_24_72 bl_int_23_72 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c73
+ bl_int_24_73 bl_int_23_73 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c74
+ bl_int_24_74 bl_int_23_74 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c75
+ bl_int_24_75 bl_int_23_75 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c76
+ bl_int_24_76 bl_int_23_76 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c77
+ bl_int_24_77 bl_int_23_77 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c78
+ bl_int_24_78 bl_int_23_78 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c79
+ bl_int_24_79 bl_int_23_79 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c80
+ bl_int_24_80 bl_int_23_80 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c81
+ bl_int_24_81 bl_int_23_81 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c82
+ bl_int_24_82 bl_int_23_82 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c83
+ bl_int_24_83 bl_int_23_83 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c84
+ bl_int_24_84 bl_int_23_84 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c85
+ bl_int_24_85 bl_int_23_85 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c86
+ bl_int_24_86 bl_int_23_86 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c87
+ bl_int_24_87 bl_int_23_87 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c88
+ bl_int_24_88 bl_int_23_88 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c89
+ bl_int_24_89 bl_int_23_89 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c90
+ bl_int_24_90 bl_int_23_90 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c91
+ bl_int_24_91 bl_int_23_91 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c92
+ bl_int_24_92 bl_int_23_92 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c93
+ bl_int_24_93 bl_int_23_93 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c94
+ bl_int_24_94 bl_int_23_94 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c95
+ bl_int_24_95 bl_int_23_95 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c96
+ bl_int_24_96 bl_int_23_96 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c97
+ bl_int_24_97 bl_int_23_97 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c98
+ bl_int_24_98 bl_int_23_98 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c99
+ bl_int_24_99 bl_int_23_99 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c100
+ bl_int_24_100 bl_int_23_100 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c101
+ bl_int_24_101 bl_int_23_101 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c102
+ bl_int_24_102 bl_int_23_102 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c103
+ bl_int_24_103 bl_int_23_103 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c104
+ bl_int_24_104 bl_int_23_104 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c105
+ bl_int_24_105 bl_int_23_105 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c106
+ bl_int_24_106 bl_int_23_106 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c107
+ bl_int_24_107 bl_int_23_107 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c108
+ bl_int_24_108 bl_int_23_108 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c109
+ bl_int_24_109 bl_int_23_109 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c110
+ bl_int_24_110 bl_int_23_110 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c111
+ bl_int_24_111 bl_int_23_111 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c112
+ bl_int_24_112 bl_int_23_112 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c113
+ bl_int_24_113 bl_int_23_113 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c114
+ bl_int_24_114 bl_int_23_114 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c115
+ bl_int_24_115 bl_int_23_115 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c116
+ bl_int_24_116 bl_int_23_116 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c117
+ bl_int_24_117 bl_int_23_117 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c118
+ bl_int_24_118 bl_int_23_118 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c119
+ bl_int_24_119 bl_int_23_119 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c120
+ bl_int_24_120 bl_int_23_120 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c121
+ bl_int_24_121 bl_int_23_121 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c122
+ bl_int_24_122 bl_int_23_122 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c123
+ bl_int_24_123 bl_int_23_123 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c124
+ bl_int_24_124 bl_int_23_124 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c125
+ bl_int_24_125 bl_int_23_125 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c126
+ bl_int_24_126 bl_int_23_126 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c127
+ bl_int_24_127 bl_int_23_127 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c128
+ bl_int_24_128 bl_int_23_128 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c129
+ bl_int_24_129 bl_int_23_129 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c130
+ bl_int_24_130 bl_int_23_130 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c131
+ bl_int_24_131 bl_int_23_131 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c132
+ bl_int_24_132 bl_int_23_132 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c133
+ bl_int_24_133 bl_int_23_133 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c134
+ bl_int_24_134 bl_int_23_134 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c135
+ bl_int_24_135 bl_int_23_135 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c136
+ bl_int_24_136 bl_int_23_136 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c137
+ bl_int_24_137 bl_int_23_137 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c138
+ bl_int_24_138 bl_int_23_138 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c139
+ bl_int_24_139 bl_int_23_139 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c140
+ bl_int_24_140 bl_int_23_140 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c141
+ bl_int_24_141 bl_int_23_141 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c142
+ bl_int_24_142 bl_int_23_142 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c143
+ bl_int_24_143 bl_int_23_143 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c144
+ bl_int_24_144 bl_int_23_144 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c145
+ bl_int_24_145 bl_int_23_145 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c146
+ bl_int_24_146 bl_int_23_146 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c147
+ bl_int_24_147 bl_int_23_147 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c148
+ bl_int_24_148 bl_int_23_148 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c149
+ bl_int_24_149 bl_int_23_149 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c150
+ bl_int_24_150 bl_int_23_150 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c151
+ bl_int_24_151 bl_int_23_151 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c152
+ bl_int_24_152 bl_int_23_152 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c153
+ bl_int_24_153 bl_int_23_153 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c154
+ bl_int_24_154 bl_int_23_154 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c155
+ bl_int_24_155 bl_int_23_155 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c156
+ bl_int_24_156 bl_int_23_156 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c157
+ bl_int_24_157 bl_int_23_157 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c158
+ bl_int_24_158 bl_int_23_158 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c159
+ bl_int_24_159 bl_int_23_159 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c160
+ bl_int_24_160 bl_int_23_160 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c161
+ bl_int_24_161 bl_int_23_161 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c162
+ bl_int_24_162 bl_int_23_162 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c163
+ bl_int_24_163 bl_int_23_163 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c164
+ bl_int_24_164 bl_int_23_164 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c165
+ bl_int_24_165 bl_int_23_165 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c166
+ bl_int_24_166 bl_int_23_166 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c167
+ bl_int_24_167 bl_int_23_167 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c168
+ bl_int_24_168 bl_int_23_168 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c169
+ bl_int_24_169 bl_int_23_169 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c170
+ bl_int_24_170 bl_int_23_170 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c171
+ bl_int_24_171 bl_int_23_171 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c172
+ bl_int_24_172 bl_int_23_172 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c173
+ bl_int_24_173 bl_int_23_173 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c174
+ bl_int_24_174 bl_int_23_174 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c175
+ bl_int_24_175 bl_int_23_175 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c176
+ bl_int_24_176 bl_int_23_176 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c177
+ bl_int_24_177 bl_int_23_177 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c178
+ bl_int_24_178 bl_int_23_178 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c179
+ bl_int_24_179 bl_int_23_179 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c180
+ bl_int_24_180 bl_int_23_180 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c181
+ bl_int_24_181 bl_int_23_181 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c182
+ bl_int_24_182 bl_int_23_182 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r24_c183
+ bl_int_24_183 bl_int_23_183 wl_0_24 gnd
+ sram_rom_base_one_cell
Xbit_r25_c0
+ bl_int_25_0 bl_int_24_0 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c1
+ bl_int_25_1 bl_int_24_1 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c2
+ bl_int_25_2 bl_int_24_2 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c3
+ bl_int_25_3 bl_int_24_3 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c4
+ bl_int_25_4 bl_int_24_4 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c5
+ bl_int_25_5 bl_int_24_5 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c6
+ bl_int_25_6 bl_int_24_6 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c7
+ bl_int_25_7 bl_int_24_7 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c8
+ bl_int_25_8 bl_int_24_8 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c9
+ bl_int_25_9 bl_int_24_9 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c10
+ bl_int_25_10 bl_int_24_10 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c11
+ bl_int_25_11 bl_int_24_11 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c12
+ bl_int_25_12 bl_int_24_12 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c13
+ bl_int_25_13 bl_int_24_13 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c14
+ bl_int_25_14 bl_int_24_14 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c15
+ bl_int_25_15 bl_int_24_15 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c16
+ bl_int_25_16 bl_int_24_16 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c17
+ bl_int_25_17 bl_int_24_17 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c18
+ bl_int_25_18 bl_int_24_18 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c19
+ bl_int_25_19 bl_int_24_19 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c20
+ bl_int_25_20 bl_int_24_20 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c21
+ bl_int_25_21 bl_int_24_21 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c22
+ bl_int_25_22 bl_int_24_22 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c23
+ bl_int_25_23 bl_int_24_23 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c24
+ bl_int_25_24 bl_int_24_24 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c25
+ bl_int_25_25 bl_int_24_25 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c26
+ bl_int_25_26 bl_int_24_26 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c27
+ bl_int_25_27 bl_int_24_27 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c28
+ bl_int_25_28 bl_int_24_28 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c29
+ bl_int_25_29 bl_int_24_29 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c30
+ bl_int_25_30 bl_int_24_30 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c31
+ bl_int_25_31 bl_int_24_31 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c32
+ bl_int_25_32 bl_int_24_32 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c33
+ bl_int_25_33 bl_int_24_33 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c34
+ bl_int_25_34 bl_int_24_34 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c35
+ bl_int_25_35 bl_int_24_35 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c36
+ bl_int_25_36 bl_int_24_36 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c37
+ bl_int_25_37 bl_int_24_37 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c38
+ bl_int_25_38 bl_int_24_38 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c39
+ bl_int_25_39 bl_int_24_39 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c40
+ bl_int_25_40 bl_int_24_40 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c41
+ bl_int_25_41 bl_int_24_41 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c42
+ bl_int_25_42 bl_int_24_42 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c43
+ bl_int_25_43 bl_int_24_43 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c44
+ bl_int_25_44 bl_int_24_44 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c45
+ bl_int_25_45 bl_int_24_45 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c46
+ bl_int_25_46 bl_int_24_46 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c47
+ bl_int_25_47 bl_int_24_47 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c48
+ bl_int_25_48 bl_int_24_48 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c49
+ bl_int_25_49 bl_int_24_49 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c50
+ bl_int_25_50 bl_int_24_50 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c51
+ bl_int_25_51 bl_int_24_51 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c52
+ bl_int_25_52 bl_int_24_52 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c53
+ bl_int_25_53 bl_int_24_53 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c54
+ bl_int_25_54 bl_int_24_54 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c55
+ bl_int_25_55 bl_int_24_55 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c56
+ bl_int_25_56 bl_int_24_56 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c57
+ bl_int_25_57 bl_int_24_57 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c58
+ bl_int_25_58 bl_int_24_58 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c59
+ bl_int_25_59 bl_int_24_59 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c60
+ bl_int_25_60 bl_int_24_60 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c61
+ bl_int_25_61 bl_int_24_61 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c62
+ bl_int_25_62 bl_int_24_62 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c63
+ bl_int_25_63 bl_int_24_63 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c64
+ bl_int_25_64 bl_int_24_64 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c65
+ bl_int_25_65 bl_int_24_65 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c66
+ bl_int_25_66 bl_int_24_66 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c67
+ bl_int_25_67 bl_int_24_67 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c68
+ bl_int_25_68 bl_int_24_68 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c69
+ bl_int_25_69 bl_int_24_69 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c70
+ bl_int_25_70 bl_int_24_70 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c71
+ bl_int_25_71 bl_int_24_71 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c72
+ bl_int_25_72 bl_int_24_72 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c73
+ bl_int_25_73 bl_int_24_73 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c74
+ bl_int_25_74 bl_int_24_74 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c75
+ bl_int_25_75 bl_int_24_75 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c76
+ bl_int_25_76 bl_int_24_76 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c77
+ bl_int_25_77 bl_int_24_77 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c78
+ bl_int_25_78 bl_int_24_78 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c79
+ bl_int_25_79 bl_int_24_79 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c80
+ bl_int_25_80 bl_int_24_80 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c81
+ bl_int_25_81 bl_int_24_81 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c82
+ bl_int_25_82 bl_int_24_82 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c83
+ bl_int_25_83 bl_int_24_83 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c84
+ bl_int_25_84 bl_int_24_84 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c85
+ bl_int_25_85 bl_int_24_85 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c86
+ bl_int_25_86 bl_int_24_86 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c87
+ bl_int_25_87 bl_int_24_87 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c88
+ bl_int_25_88 bl_int_24_88 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c89
+ bl_int_25_89 bl_int_24_89 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c90
+ bl_int_25_90 bl_int_24_90 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c91
+ bl_int_25_91 bl_int_24_91 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c92
+ bl_int_25_92 bl_int_24_92 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c93
+ bl_int_25_93 bl_int_24_93 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c94
+ bl_int_25_94 bl_int_24_94 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c95
+ bl_int_25_95 bl_int_24_95 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c96
+ bl_int_25_96 bl_int_24_96 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c97
+ bl_int_25_97 bl_int_24_97 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c98
+ bl_int_25_98 bl_int_24_98 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c99
+ bl_int_25_99 bl_int_24_99 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c100
+ bl_int_25_100 bl_int_24_100 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c101
+ bl_int_25_101 bl_int_24_101 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c102
+ bl_int_25_102 bl_int_24_102 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c103
+ bl_int_25_103 bl_int_24_103 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c104
+ bl_int_25_104 bl_int_24_104 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c105
+ bl_int_25_105 bl_int_24_105 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c106
+ bl_int_25_106 bl_int_24_106 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c107
+ bl_int_25_107 bl_int_24_107 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c108
+ bl_int_25_108 bl_int_24_108 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c109
+ bl_int_25_109 bl_int_24_109 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c110
+ bl_int_25_110 bl_int_24_110 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c111
+ bl_int_25_111 bl_int_24_111 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c112
+ bl_int_25_112 bl_int_24_112 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c113
+ bl_int_25_113 bl_int_24_113 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c114
+ bl_int_25_114 bl_int_24_114 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c115
+ bl_int_25_115 bl_int_24_115 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c116
+ bl_int_25_116 bl_int_24_116 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c117
+ bl_int_25_117 bl_int_24_117 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c118
+ bl_int_25_118 bl_int_24_118 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c119
+ bl_int_25_119 bl_int_24_119 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c120
+ bl_int_25_120 bl_int_24_120 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c121
+ bl_int_25_121 bl_int_24_121 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c122
+ bl_int_25_122 bl_int_24_122 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c123
+ bl_int_25_123 bl_int_24_123 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c124
+ bl_int_25_124 bl_int_24_124 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c125
+ bl_int_25_125 bl_int_24_125 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c126
+ bl_int_25_126 bl_int_24_126 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c127
+ bl_int_25_127 bl_int_24_127 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c128
+ bl_int_25_128 bl_int_24_128 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c129
+ bl_int_25_129 bl_int_24_129 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c130
+ bl_int_25_130 bl_int_24_130 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c131
+ bl_int_25_131 bl_int_24_131 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c132
+ bl_int_25_132 bl_int_24_132 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c133
+ bl_int_25_133 bl_int_24_133 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c134
+ bl_int_25_134 bl_int_24_134 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c135
+ bl_int_25_135 bl_int_24_135 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c136
+ bl_int_25_136 bl_int_24_136 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c137
+ bl_int_25_137 bl_int_24_137 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c138
+ bl_int_25_138 bl_int_24_138 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c139
+ bl_int_25_139 bl_int_24_139 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c140
+ bl_int_25_140 bl_int_24_140 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c141
+ bl_int_25_141 bl_int_24_141 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c142
+ bl_int_25_142 bl_int_24_142 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c143
+ bl_int_25_143 bl_int_24_143 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c144
+ bl_int_25_144 bl_int_24_144 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c145
+ bl_int_25_145 bl_int_24_145 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c146
+ bl_int_25_146 bl_int_24_146 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c147
+ bl_int_25_147 bl_int_24_147 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c148
+ bl_int_25_148 bl_int_24_148 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c149
+ bl_int_25_149 bl_int_24_149 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c150
+ bl_int_25_150 bl_int_24_150 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c151
+ bl_int_25_151 bl_int_24_151 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c152
+ bl_int_25_152 bl_int_24_152 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c153
+ bl_int_25_153 bl_int_24_153 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c154
+ bl_int_25_154 bl_int_24_154 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c155
+ bl_int_25_155 bl_int_24_155 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c156
+ bl_int_25_156 bl_int_24_156 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c157
+ bl_int_25_157 bl_int_24_157 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c158
+ bl_int_25_158 bl_int_24_158 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c159
+ bl_int_25_159 bl_int_24_159 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c160
+ bl_int_25_160 bl_int_24_160 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c161
+ bl_int_25_161 bl_int_24_161 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c162
+ bl_int_25_162 bl_int_24_162 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c163
+ bl_int_25_163 bl_int_24_163 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c164
+ bl_int_25_164 bl_int_24_164 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c165
+ bl_int_25_165 bl_int_24_165 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c166
+ bl_int_25_166 bl_int_24_166 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c167
+ bl_int_25_167 bl_int_24_167 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c168
+ bl_int_25_168 bl_int_24_168 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c169
+ bl_int_25_169 bl_int_24_169 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c170
+ bl_int_25_170 bl_int_24_170 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c171
+ bl_int_25_171 bl_int_24_171 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c172
+ bl_int_25_172 bl_int_24_172 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c173
+ bl_int_25_173 bl_int_24_173 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c174
+ bl_int_25_174 bl_int_24_174 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c175
+ bl_int_25_175 bl_int_24_175 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c176
+ bl_int_25_176 bl_int_24_176 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c177
+ bl_int_25_177 bl_int_24_177 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c178
+ bl_int_25_178 bl_int_24_178 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c179
+ bl_int_25_179 bl_int_24_179 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c180
+ bl_int_25_180 bl_int_24_180 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c181
+ bl_int_25_181 bl_int_24_181 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c182
+ bl_int_25_182 bl_int_24_182 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r25_c183
+ bl_int_25_183 bl_int_24_183 wl_0_25 gnd
+ sram_rom_base_one_cell
Xbit_r26_c0
+ bl_int_26_0 bl_int_25_0 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c1
+ bl_int_26_1 bl_int_25_1 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c2
+ bl_int_26_2 bl_int_25_2 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c3
+ bl_int_26_3 bl_int_25_3 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c4
+ bl_int_26_4 bl_int_25_4 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c5
+ bl_int_26_5 bl_int_25_5 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c6
+ bl_int_26_6 bl_int_25_6 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c7
+ bl_int_26_7 bl_int_25_7 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c8
+ bl_int_26_8 bl_int_25_8 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c9
+ bl_int_26_9 bl_int_25_9 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c10
+ bl_int_26_10 bl_int_25_10 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c11
+ bl_int_26_11 bl_int_25_11 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c12
+ bl_int_26_12 bl_int_25_12 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c13
+ bl_int_26_13 bl_int_25_13 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c14
+ bl_int_26_14 bl_int_25_14 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c15
+ bl_int_26_15 bl_int_25_15 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c16
+ bl_int_26_16 bl_int_25_16 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c17
+ bl_int_26_17 bl_int_25_17 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c18
+ bl_int_26_18 bl_int_25_18 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c19
+ bl_int_26_19 bl_int_25_19 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c20
+ bl_int_26_20 bl_int_25_20 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c21
+ bl_int_26_21 bl_int_25_21 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c22
+ bl_int_26_22 bl_int_25_22 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c23
+ bl_int_26_23 bl_int_25_23 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c24
+ bl_int_26_24 bl_int_25_24 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c25
+ bl_int_26_25 bl_int_25_25 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c26
+ bl_int_26_26 bl_int_25_26 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c27
+ bl_int_26_27 bl_int_25_27 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c28
+ bl_int_26_28 bl_int_25_28 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c29
+ bl_int_26_29 bl_int_25_29 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c30
+ bl_int_26_30 bl_int_25_30 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c31
+ bl_int_26_31 bl_int_25_31 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c32
+ bl_int_26_32 bl_int_25_32 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c33
+ bl_int_26_33 bl_int_25_33 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c34
+ bl_int_26_34 bl_int_25_34 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c35
+ bl_int_26_35 bl_int_25_35 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c36
+ bl_int_26_36 bl_int_25_36 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c37
+ bl_int_26_37 bl_int_25_37 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c38
+ bl_int_26_38 bl_int_25_38 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c39
+ bl_int_26_39 bl_int_25_39 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c40
+ bl_int_26_40 bl_int_25_40 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c41
+ bl_int_26_41 bl_int_25_41 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c42
+ bl_int_26_42 bl_int_25_42 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c43
+ bl_int_26_43 bl_int_25_43 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c44
+ bl_int_26_44 bl_int_25_44 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c45
+ bl_int_26_45 bl_int_25_45 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c46
+ bl_int_26_46 bl_int_25_46 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c47
+ bl_int_26_47 bl_int_25_47 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c48
+ bl_int_26_48 bl_int_25_48 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c49
+ bl_int_26_49 bl_int_25_49 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c50
+ bl_int_26_50 bl_int_25_50 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c51
+ bl_int_26_51 bl_int_25_51 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c52
+ bl_int_26_52 bl_int_25_52 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c53
+ bl_int_26_53 bl_int_25_53 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c54
+ bl_int_26_54 bl_int_25_54 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c55
+ bl_int_26_55 bl_int_25_55 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c56
+ bl_int_26_56 bl_int_25_56 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c57
+ bl_int_26_57 bl_int_25_57 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c58
+ bl_int_26_58 bl_int_25_58 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c59
+ bl_int_26_59 bl_int_25_59 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c60
+ bl_int_26_60 bl_int_25_60 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c61
+ bl_int_26_61 bl_int_25_61 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c62
+ bl_int_26_62 bl_int_25_62 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c63
+ bl_int_26_63 bl_int_25_63 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c64
+ bl_int_26_64 bl_int_25_64 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c65
+ bl_int_26_65 bl_int_25_65 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c66
+ bl_int_26_66 bl_int_25_66 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c67
+ bl_int_26_67 bl_int_25_67 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c68
+ bl_int_26_68 bl_int_25_68 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c69
+ bl_int_26_69 bl_int_25_69 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c70
+ bl_int_26_70 bl_int_25_70 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c71
+ bl_int_26_71 bl_int_25_71 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c72
+ bl_int_26_72 bl_int_25_72 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c73
+ bl_int_26_73 bl_int_25_73 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c74
+ bl_int_26_74 bl_int_25_74 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c75
+ bl_int_26_75 bl_int_25_75 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c76
+ bl_int_26_76 bl_int_25_76 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c77
+ bl_int_26_77 bl_int_25_77 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c78
+ bl_int_26_78 bl_int_25_78 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c79
+ bl_int_26_79 bl_int_25_79 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c80
+ bl_int_26_80 bl_int_25_80 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c81
+ bl_int_26_81 bl_int_25_81 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c82
+ bl_int_26_82 bl_int_25_82 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c83
+ bl_int_26_83 bl_int_25_83 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c84
+ bl_int_26_84 bl_int_25_84 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c85
+ bl_int_26_85 bl_int_25_85 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c86
+ bl_int_26_86 bl_int_25_86 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c87
+ bl_int_26_87 bl_int_25_87 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c88
+ bl_int_26_88 bl_int_25_88 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c89
+ bl_int_26_89 bl_int_25_89 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c90
+ bl_int_26_90 bl_int_25_90 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c91
+ bl_int_26_91 bl_int_25_91 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c92
+ bl_int_26_92 bl_int_25_92 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c93
+ bl_int_26_93 bl_int_25_93 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c94
+ bl_int_26_94 bl_int_25_94 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c95
+ bl_int_26_95 bl_int_25_95 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c96
+ bl_int_26_96 bl_int_25_96 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c97
+ bl_int_26_97 bl_int_25_97 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c98
+ bl_int_26_98 bl_int_25_98 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c99
+ bl_int_26_99 bl_int_25_99 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c100
+ bl_int_26_100 bl_int_25_100 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c101
+ bl_int_26_101 bl_int_25_101 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c102
+ bl_int_26_102 bl_int_25_102 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c103
+ bl_int_26_103 bl_int_25_103 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c104
+ bl_int_26_104 bl_int_25_104 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c105
+ bl_int_26_105 bl_int_25_105 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c106
+ bl_int_26_106 bl_int_25_106 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c107
+ bl_int_26_107 bl_int_25_107 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c108
+ bl_int_26_108 bl_int_25_108 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c109
+ bl_int_26_109 bl_int_25_109 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c110
+ bl_int_26_110 bl_int_25_110 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c111
+ bl_int_26_111 bl_int_25_111 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c112
+ bl_int_26_112 bl_int_25_112 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c113
+ bl_int_26_113 bl_int_25_113 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c114
+ bl_int_26_114 bl_int_25_114 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c115
+ bl_int_26_115 bl_int_25_115 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c116
+ bl_int_26_116 bl_int_25_116 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c117
+ bl_int_26_117 bl_int_25_117 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c118
+ bl_int_26_118 bl_int_25_118 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c119
+ bl_int_26_119 bl_int_25_119 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c120
+ bl_int_26_120 bl_int_25_120 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c121
+ bl_int_26_121 bl_int_25_121 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c122
+ bl_int_26_122 bl_int_25_122 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c123
+ bl_int_26_123 bl_int_25_123 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c124
+ bl_int_26_124 bl_int_25_124 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c125
+ bl_int_26_125 bl_int_25_125 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c126
+ bl_int_26_126 bl_int_25_126 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c127
+ bl_int_26_127 bl_int_25_127 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c128
+ bl_int_26_128 bl_int_25_128 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c129
+ bl_int_26_129 bl_int_25_129 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c130
+ bl_int_26_130 bl_int_25_130 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c131
+ bl_int_26_131 bl_int_25_131 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c132
+ bl_int_26_132 bl_int_25_132 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c133
+ bl_int_26_133 bl_int_25_133 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c134
+ bl_int_26_134 bl_int_25_134 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c135
+ bl_int_26_135 bl_int_25_135 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c136
+ bl_int_26_136 bl_int_25_136 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c137
+ bl_int_26_137 bl_int_25_137 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c138
+ bl_int_26_138 bl_int_25_138 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c139
+ bl_int_26_139 bl_int_25_139 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c140
+ bl_int_26_140 bl_int_25_140 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c141
+ bl_int_26_141 bl_int_25_141 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c142
+ bl_int_26_142 bl_int_25_142 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c143
+ bl_int_26_143 bl_int_25_143 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c144
+ bl_int_26_144 bl_int_25_144 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c145
+ bl_int_26_145 bl_int_25_145 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c146
+ bl_int_26_146 bl_int_25_146 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c147
+ bl_int_26_147 bl_int_25_147 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c148
+ bl_int_26_148 bl_int_25_148 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c149
+ bl_int_26_149 bl_int_25_149 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c150
+ bl_int_26_150 bl_int_25_150 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c151
+ bl_int_26_151 bl_int_25_151 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c152
+ bl_int_26_152 bl_int_25_152 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c153
+ bl_int_26_153 bl_int_25_153 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c154
+ bl_int_26_154 bl_int_25_154 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c155
+ bl_int_26_155 bl_int_25_155 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c156
+ bl_int_26_156 bl_int_25_156 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c157
+ bl_int_26_157 bl_int_25_157 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c158
+ bl_int_26_158 bl_int_25_158 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c159
+ bl_int_26_159 bl_int_25_159 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c160
+ bl_int_26_160 bl_int_25_160 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c161
+ bl_int_26_161 bl_int_25_161 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c162
+ bl_int_26_162 bl_int_25_162 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c163
+ bl_int_26_163 bl_int_25_163 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c164
+ bl_int_26_164 bl_int_25_164 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c165
+ bl_int_26_165 bl_int_25_165 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c166
+ bl_int_26_166 bl_int_25_166 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c167
+ bl_int_26_167 bl_int_25_167 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c168
+ bl_int_26_168 bl_int_25_168 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c169
+ bl_int_26_169 bl_int_25_169 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c170
+ bl_int_26_170 bl_int_25_170 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c171
+ bl_int_26_171 bl_int_25_171 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c172
+ bl_int_26_172 bl_int_25_172 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c173
+ bl_int_26_173 bl_int_25_173 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c174
+ bl_int_26_174 bl_int_25_174 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c175
+ bl_int_26_175 bl_int_25_175 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c176
+ bl_int_26_176 bl_int_25_176 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c177
+ bl_int_26_177 bl_int_25_177 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c178
+ bl_int_26_178 bl_int_25_178 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c179
+ bl_int_26_179 bl_int_25_179 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c180
+ bl_int_26_180 bl_int_25_180 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c181
+ bl_int_26_181 bl_int_25_181 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c182
+ bl_int_26_182 bl_int_25_182 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r26_c183
+ bl_int_26_183 bl_int_25_183 wl_0_26 gnd
+ sram_rom_base_one_cell
Xbit_r27_c0
+ bl_int_27_0 bl_int_26_0 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c1
+ bl_int_27_1 bl_int_26_1 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c2
+ bl_int_27_2 bl_int_26_2 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c3
+ bl_int_27_3 bl_int_26_3 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c4
+ bl_int_27_4 bl_int_26_4 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c5
+ bl_int_27_5 bl_int_26_5 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c6
+ bl_int_27_6 bl_int_26_6 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c7
+ bl_int_27_7 bl_int_26_7 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c8
+ bl_int_27_8 bl_int_26_8 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c9
+ bl_int_27_9 bl_int_26_9 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c10
+ bl_int_27_10 bl_int_26_10 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c11
+ bl_int_27_11 bl_int_26_11 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c12
+ bl_int_27_12 bl_int_26_12 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c13
+ bl_int_27_13 bl_int_26_13 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c14
+ bl_int_27_14 bl_int_26_14 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c15
+ bl_int_27_15 bl_int_26_15 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c16
+ bl_int_27_16 bl_int_26_16 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c17
+ bl_int_27_17 bl_int_26_17 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c18
+ bl_int_27_18 bl_int_26_18 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c19
+ bl_int_27_19 bl_int_26_19 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c20
+ bl_int_27_20 bl_int_26_20 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c21
+ bl_int_27_21 bl_int_26_21 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c22
+ bl_int_27_22 bl_int_26_22 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c23
+ bl_int_27_23 bl_int_26_23 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c24
+ bl_int_27_24 bl_int_26_24 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c25
+ bl_int_27_25 bl_int_26_25 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c26
+ bl_int_27_26 bl_int_26_26 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c27
+ bl_int_27_27 bl_int_26_27 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c28
+ bl_int_27_28 bl_int_26_28 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c29
+ bl_int_27_29 bl_int_26_29 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c30
+ bl_int_27_30 bl_int_26_30 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c31
+ bl_int_27_31 bl_int_26_31 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c32
+ bl_int_27_32 bl_int_26_32 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c33
+ bl_int_27_33 bl_int_26_33 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c34
+ bl_int_27_34 bl_int_26_34 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c35
+ bl_int_27_35 bl_int_26_35 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c36
+ bl_int_27_36 bl_int_26_36 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c37
+ bl_int_27_37 bl_int_26_37 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c38
+ bl_int_27_38 bl_int_26_38 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c39
+ bl_int_27_39 bl_int_26_39 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c40
+ bl_int_27_40 bl_int_26_40 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c41
+ bl_int_27_41 bl_int_26_41 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c42
+ bl_int_27_42 bl_int_26_42 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c43
+ bl_int_27_43 bl_int_26_43 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c44
+ bl_int_27_44 bl_int_26_44 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c45
+ bl_int_27_45 bl_int_26_45 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c46
+ bl_int_27_46 bl_int_26_46 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c47
+ bl_int_27_47 bl_int_26_47 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c48
+ bl_int_27_48 bl_int_26_48 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c49
+ bl_int_27_49 bl_int_26_49 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c50
+ bl_int_27_50 bl_int_26_50 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c51
+ bl_int_27_51 bl_int_26_51 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c52
+ bl_int_27_52 bl_int_26_52 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c53
+ bl_int_27_53 bl_int_26_53 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c54
+ bl_int_27_54 bl_int_26_54 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c55
+ bl_int_27_55 bl_int_26_55 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c56
+ bl_int_27_56 bl_int_26_56 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c57
+ bl_int_27_57 bl_int_26_57 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c58
+ bl_int_27_58 bl_int_26_58 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c59
+ bl_int_27_59 bl_int_26_59 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c60
+ bl_int_27_60 bl_int_26_60 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c61
+ bl_int_27_61 bl_int_26_61 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c62
+ bl_int_27_62 bl_int_26_62 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c63
+ bl_int_27_63 bl_int_26_63 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c64
+ bl_int_27_64 bl_int_26_64 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c65
+ bl_int_27_65 bl_int_26_65 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c66
+ bl_int_27_66 bl_int_26_66 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c67
+ bl_int_27_67 bl_int_26_67 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c68
+ bl_int_27_68 bl_int_26_68 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c69
+ bl_int_27_69 bl_int_26_69 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c70
+ bl_int_27_70 bl_int_26_70 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c71
+ bl_int_27_71 bl_int_26_71 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c72
+ bl_int_27_72 bl_int_26_72 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c73
+ bl_int_27_73 bl_int_26_73 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c74
+ bl_int_27_74 bl_int_26_74 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c75
+ bl_int_27_75 bl_int_26_75 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c76
+ bl_int_27_76 bl_int_26_76 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c77
+ bl_int_27_77 bl_int_26_77 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c78
+ bl_int_27_78 bl_int_26_78 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c79
+ bl_int_27_79 bl_int_26_79 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c80
+ bl_int_27_80 bl_int_26_80 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c81
+ bl_int_27_81 bl_int_26_81 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c82
+ bl_int_27_82 bl_int_26_82 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c83
+ bl_int_27_83 bl_int_26_83 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c84
+ bl_int_27_84 bl_int_26_84 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c85
+ bl_int_27_85 bl_int_26_85 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c86
+ bl_int_27_86 bl_int_26_86 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c87
+ bl_int_27_87 bl_int_26_87 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c88
+ bl_int_27_88 bl_int_26_88 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c89
+ bl_int_27_89 bl_int_26_89 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c90
+ bl_int_27_90 bl_int_26_90 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c91
+ bl_int_27_91 bl_int_26_91 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c92
+ bl_int_27_92 bl_int_26_92 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c93
+ bl_int_27_93 bl_int_26_93 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c94
+ bl_int_27_94 bl_int_26_94 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c95
+ bl_int_27_95 bl_int_26_95 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c96
+ bl_int_27_96 bl_int_26_96 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c97
+ bl_int_27_97 bl_int_26_97 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c98
+ bl_int_27_98 bl_int_26_98 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c99
+ bl_int_27_99 bl_int_26_99 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c100
+ bl_int_27_100 bl_int_26_100 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c101
+ bl_int_27_101 bl_int_26_101 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c102
+ bl_int_27_102 bl_int_26_102 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c103
+ bl_int_27_103 bl_int_26_103 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c104
+ bl_int_27_104 bl_int_26_104 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c105
+ bl_int_27_105 bl_int_26_105 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c106
+ bl_int_27_106 bl_int_26_106 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c107
+ bl_int_27_107 bl_int_26_107 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c108
+ bl_int_27_108 bl_int_26_108 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c109
+ bl_int_27_109 bl_int_26_109 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c110
+ bl_int_27_110 bl_int_26_110 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c111
+ bl_int_27_111 bl_int_26_111 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c112
+ bl_int_27_112 bl_int_26_112 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c113
+ bl_int_27_113 bl_int_26_113 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c114
+ bl_int_27_114 bl_int_26_114 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c115
+ bl_int_27_115 bl_int_26_115 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c116
+ bl_int_27_116 bl_int_26_116 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c117
+ bl_int_27_117 bl_int_26_117 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c118
+ bl_int_27_118 bl_int_26_118 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c119
+ bl_int_27_119 bl_int_26_119 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c120
+ bl_int_27_120 bl_int_26_120 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c121
+ bl_int_27_121 bl_int_26_121 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c122
+ bl_int_27_122 bl_int_26_122 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c123
+ bl_int_27_123 bl_int_26_123 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c124
+ bl_int_27_124 bl_int_26_124 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c125
+ bl_int_27_125 bl_int_26_125 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c126
+ bl_int_27_126 bl_int_26_126 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c127
+ bl_int_27_127 bl_int_26_127 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c128
+ bl_int_27_128 bl_int_26_128 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c129
+ bl_int_27_129 bl_int_26_129 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c130
+ bl_int_27_130 bl_int_26_130 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c131
+ bl_int_27_131 bl_int_26_131 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c132
+ bl_int_27_132 bl_int_26_132 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c133
+ bl_int_27_133 bl_int_26_133 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c134
+ bl_int_27_134 bl_int_26_134 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c135
+ bl_int_27_135 bl_int_26_135 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c136
+ bl_int_27_136 bl_int_26_136 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c137
+ bl_int_27_137 bl_int_26_137 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c138
+ bl_int_27_138 bl_int_26_138 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c139
+ bl_int_27_139 bl_int_26_139 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c140
+ bl_int_27_140 bl_int_26_140 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c141
+ bl_int_27_141 bl_int_26_141 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c142
+ bl_int_27_142 bl_int_26_142 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c143
+ bl_int_27_143 bl_int_26_143 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c144
+ bl_int_27_144 bl_int_26_144 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c145
+ bl_int_27_145 bl_int_26_145 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c146
+ bl_int_27_146 bl_int_26_146 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c147
+ bl_int_27_147 bl_int_26_147 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c148
+ bl_int_27_148 bl_int_26_148 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c149
+ bl_int_27_149 bl_int_26_149 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c150
+ bl_int_27_150 bl_int_26_150 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c151
+ bl_int_27_151 bl_int_26_151 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c152
+ bl_int_27_152 bl_int_26_152 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c153
+ bl_int_27_153 bl_int_26_153 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c154
+ bl_int_27_154 bl_int_26_154 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c155
+ bl_int_27_155 bl_int_26_155 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c156
+ bl_int_27_156 bl_int_26_156 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c157
+ bl_int_27_157 bl_int_26_157 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c158
+ bl_int_27_158 bl_int_26_158 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c159
+ bl_int_27_159 bl_int_26_159 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c160
+ bl_int_27_160 bl_int_26_160 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c161
+ bl_int_27_161 bl_int_26_161 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c162
+ bl_int_27_162 bl_int_26_162 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c163
+ bl_int_27_163 bl_int_26_163 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c164
+ bl_int_27_164 bl_int_26_164 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c165
+ bl_int_27_165 bl_int_26_165 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c166
+ bl_int_27_166 bl_int_26_166 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c167
+ bl_int_27_167 bl_int_26_167 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c168
+ bl_int_27_168 bl_int_26_168 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c169
+ bl_int_27_169 bl_int_26_169 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c170
+ bl_int_27_170 bl_int_26_170 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c171
+ bl_int_27_171 bl_int_26_171 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c172
+ bl_int_27_172 bl_int_26_172 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c173
+ bl_int_27_173 bl_int_26_173 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c174
+ bl_int_27_174 bl_int_26_174 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c175
+ bl_int_27_175 bl_int_26_175 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c176
+ bl_int_27_176 bl_int_26_176 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c177
+ bl_int_27_177 bl_int_26_177 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c178
+ bl_int_27_178 bl_int_26_178 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c179
+ bl_int_27_179 bl_int_26_179 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c180
+ bl_int_27_180 bl_int_26_180 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c181
+ bl_int_27_181 bl_int_26_181 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c182
+ bl_int_27_182 bl_int_26_182 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r27_c183
+ bl_int_27_183 bl_int_26_183 wl_0_27 gnd
+ sram_rom_base_one_cell
Xbit_r28_c0
+ bl_int_28_0 bl_int_27_0 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c1
+ bl_int_28_1 bl_int_27_1 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c2
+ bl_int_28_2 bl_int_27_2 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c3
+ bl_int_28_3 bl_int_27_3 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c4
+ bl_int_28_4 bl_int_27_4 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c5
+ bl_int_28_5 bl_int_27_5 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c6
+ bl_int_28_6 bl_int_27_6 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c7
+ bl_int_28_7 bl_int_27_7 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c8
+ bl_int_28_8 bl_int_27_8 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c9
+ bl_int_28_9 bl_int_27_9 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c10
+ bl_int_28_10 bl_int_27_10 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c11
+ bl_int_28_11 bl_int_27_11 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c12
+ bl_int_28_12 bl_int_27_12 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c13
+ bl_int_28_13 bl_int_27_13 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c14
+ bl_int_28_14 bl_int_27_14 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c15
+ bl_int_28_15 bl_int_27_15 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c16
+ bl_int_28_16 bl_int_27_16 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c17
+ bl_int_28_17 bl_int_27_17 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c18
+ bl_int_28_18 bl_int_27_18 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c19
+ bl_int_28_19 bl_int_27_19 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c20
+ bl_int_28_20 bl_int_27_20 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c21
+ bl_int_28_21 bl_int_27_21 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c22
+ bl_int_28_22 bl_int_27_22 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c23
+ bl_int_28_23 bl_int_27_23 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c24
+ bl_int_28_24 bl_int_27_24 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c25
+ bl_int_28_25 bl_int_27_25 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c26
+ bl_int_28_26 bl_int_27_26 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c27
+ bl_int_28_27 bl_int_27_27 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c28
+ bl_int_28_28 bl_int_27_28 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c29
+ bl_int_28_29 bl_int_27_29 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c30
+ bl_int_28_30 bl_int_27_30 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c31
+ bl_int_28_31 bl_int_27_31 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c32
+ bl_int_28_32 bl_int_27_32 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c33
+ bl_int_28_33 bl_int_27_33 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c34
+ bl_int_28_34 bl_int_27_34 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c35
+ bl_int_28_35 bl_int_27_35 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c36
+ bl_int_28_36 bl_int_27_36 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c37
+ bl_int_28_37 bl_int_27_37 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c38
+ bl_int_28_38 bl_int_27_38 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c39
+ bl_int_28_39 bl_int_27_39 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c40
+ bl_int_28_40 bl_int_27_40 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c41
+ bl_int_28_41 bl_int_27_41 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c42
+ bl_int_28_42 bl_int_27_42 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c43
+ bl_int_28_43 bl_int_27_43 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c44
+ bl_int_28_44 bl_int_27_44 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c45
+ bl_int_28_45 bl_int_27_45 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c46
+ bl_int_28_46 bl_int_27_46 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c47
+ bl_int_28_47 bl_int_27_47 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c48
+ bl_int_28_48 bl_int_27_48 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c49
+ bl_int_28_49 bl_int_27_49 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c50
+ bl_int_28_50 bl_int_27_50 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c51
+ bl_int_28_51 bl_int_27_51 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c52
+ bl_int_28_52 bl_int_27_52 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c53
+ bl_int_28_53 bl_int_27_53 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c54
+ bl_int_28_54 bl_int_27_54 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c55
+ bl_int_28_55 bl_int_27_55 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c56
+ bl_int_28_56 bl_int_27_56 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c57
+ bl_int_28_57 bl_int_27_57 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c58
+ bl_int_28_58 bl_int_27_58 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c59
+ bl_int_28_59 bl_int_27_59 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c60
+ bl_int_28_60 bl_int_27_60 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c61
+ bl_int_28_61 bl_int_27_61 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c62
+ bl_int_28_62 bl_int_27_62 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c63
+ bl_int_28_63 bl_int_27_63 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c64
+ bl_int_28_64 bl_int_27_64 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c65
+ bl_int_28_65 bl_int_27_65 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c66
+ bl_int_28_66 bl_int_27_66 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c67
+ bl_int_28_67 bl_int_27_67 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c68
+ bl_int_28_68 bl_int_27_68 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c69
+ bl_int_28_69 bl_int_27_69 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c70
+ bl_int_28_70 bl_int_27_70 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c71
+ bl_int_28_71 bl_int_27_71 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c72
+ bl_int_28_72 bl_int_27_72 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c73
+ bl_int_28_73 bl_int_27_73 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c74
+ bl_int_28_74 bl_int_27_74 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c75
+ bl_int_28_75 bl_int_27_75 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c76
+ bl_int_28_76 bl_int_27_76 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c77
+ bl_int_28_77 bl_int_27_77 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c78
+ bl_int_28_78 bl_int_27_78 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c79
+ bl_int_28_79 bl_int_27_79 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c80
+ bl_int_28_80 bl_int_27_80 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c81
+ bl_int_28_81 bl_int_27_81 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c82
+ bl_int_28_82 bl_int_27_82 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c83
+ bl_int_28_83 bl_int_27_83 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c84
+ bl_int_28_84 bl_int_27_84 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c85
+ bl_int_28_85 bl_int_27_85 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c86
+ bl_int_28_86 bl_int_27_86 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c87
+ bl_int_28_87 bl_int_27_87 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c88
+ bl_int_28_88 bl_int_27_88 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c89
+ bl_int_28_89 bl_int_27_89 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c90
+ bl_int_28_90 bl_int_27_90 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c91
+ bl_int_28_91 bl_int_27_91 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c92
+ bl_int_28_92 bl_int_27_92 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c93
+ bl_int_28_93 bl_int_27_93 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c94
+ bl_int_28_94 bl_int_27_94 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c95
+ bl_int_28_95 bl_int_27_95 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c96
+ bl_int_28_96 bl_int_27_96 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c97
+ bl_int_28_97 bl_int_27_97 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c98
+ bl_int_28_98 bl_int_27_98 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c99
+ bl_int_28_99 bl_int_27_99 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c100
+ bl_int_28_100 bl_int_27_100 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c101
+ bl_int_28_101 bl_int_27_101 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c102
+ bl_int_28_102 bl_int_27_102 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c103
+ bl_int_28_103 bl_int_27_103 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c104
+ bl_int_28_104 bl_int_27_104 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c105
+ bl_int_28_105 bl_int_27_105 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c106
+ bl_int_28_106 bl_int_27_106 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c107
+ bl_int_28_107 bl_int_27_107 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c108
+ bl_int_28_108 bl_int_27_108 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c109
+ bl_int_28_109 bl_int_27_109 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c110
+ bl_int_28_110 bl_int_27_110 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c111
+ bl_int_28_111 bl_int_27_111 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c112
+ bl_int_28_112 bl_int_27_112 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c113
+ bl_int_28_113 bl_int_27_113 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c114
+ bl_int_28_114 bl_int_27_114 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c115
+ bl_int_28_115 bl_int_27_115 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c116
+ bl_int_28_116 bl_int_27_116 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c117
+ bl_int_28_117 bl_int_27_117 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c118
+ bl_int_28_118 bl_int_27_118 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c119
+ bl_int_28_119 bl_int_27_119 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c120
+ bl_int_28_120 bl_int_27_120 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c121
+ bl_int_28_121 bl_int_27_121 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c122
+ bl_int_28_122 bl_int_27_122 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c123
+ bl_int_28_123 bl_int_27_123 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c124
+ bl_int_28_124 bl_int_27_124 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c125
+ bl_int_28_125 bl_int_27_125 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c126
+ bl_int_28_126 bl_int_27_126 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c127
+ bl_int_28_127 bl_int_27_127 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c128
+ bl_int_28_128 bl_int_27_128 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c129
+ bl_int_28_129 bl_int_27_129 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c130
+ bl_int_28_130 bl_int_27_130 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c131
+ bl_int_28_131 bl_int_27_131 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c132
+ bl_int_28_132 bl_int_27_132 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c133
+ bl_int_28_133 bl_int_27_133 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c134
+ bl_int_28_134 bl_int_27_134 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c135
+ bl_int_28_135 bl_int_27_135 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c136
+ bl_int_28_136 bl_int_27_136 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c137
+ bl_int_28_137 bl_int_27_137 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c138
+ bl_int_28_138 bl_int_27_138 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c139
+ bl_int_28_139 bl_int_27_139 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c140
+ bl_int_28_140 bl_int_27_140 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c141
+ bl_int_28_141 bl_int_27_141 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c142
+ bl_int_28_142 bl_int_27_142 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c143
+ bl_int_28_143 bl_int_27_143 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c144
+ bl_int_28_144 bl_int_27_144 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c145
+ bl_int_28_145 bl_int_27_145 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c146
+ bl_int_28_146 bl_int_27_146 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c147
+ bl_int_28_147 bl_int_27_147 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c148
+ bl_int_28_148 bl_int_27_148 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c149
+ bl_int_28_149 bl_int_27_149 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c150
+ bl_int_28_150 bl_int_27_150 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c151
+ bl_int_28_151 bl_int_27_151 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c152
+ bl_int_28_152 bl_int_27_152 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c153
+ bl_int_28_153 bl_int_27_153 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c154
+ bl_int_28_154 bl_int_27_154 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c155
+ bl_int_28_155 bl_int_27_155 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c156
+ bl_int_28_156 bl_int_27_156 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c157
+ bl_int_28_157 bl_int_27_157 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c158
+ bl_int_28_158 bl_int_27_158 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c159
+ bl_int_28_159 bl_int_27_159 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c160
+ bl_int_28_160 bl_int_27_160 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c161
+ bl_int_28_161 bl_int_27_161 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c162
+ bl_int_28_162 bl_int_27_162 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c163
+ bl_int_28_163 bl_int_27_163 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c164
+ bl_int_28_164 bl_int_27_164 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c165
+ bl_int_28_165 bl_int_27_165 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c166
+ bl_int_28_166 bl_int_27_166 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c167
+ bl_int_28_167 bl_int_27_167 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c168
+ bl_int_28_168 bl_int_27_168 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c169
+ bl_int_28_169 bl_int_27_169 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c170
+ bl_int_28_170 bl_int_27_170 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c171
+ bl_int_28_171 bl_int_27_171 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c172
+ bl_int_28_172 bl_int_27_172 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c173
+ bl_int_28_173 bl_int_27_173 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c174
+ bl_int_28_174 bl_int_27_174 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c175
+ bl_int_28_175 bl_int_27_175 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c176
+ bl_int_28_176 bl_int_27_176 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c177
+ bl_int_28_177 bl_int_27_177 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c178
+ bl_int_28_178 bl_int_27_178 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c179
+ bl_int_28_179 bl_int_27_179 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c180
+ bl_int_28_180 bl_int_27_180 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c181
+ bl_int_28_181 bl_int_27_181 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c182
+ bl_int_28_182 bl_int_27_182 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r28_c183
+ bl_int_28_183 bl_int_27_183 wl_0_28 gnd
+ sram_rom_base_one_cell
Xbit_r29_c0
+ bl_int_29_0 bl_int_28_0 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c1
+ bl_int_29_1 bl_int_28_1 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c2
+ bl_int_29_2 bl_int_28_2 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c3
+ bl_int_29_3 bl_int_28_3 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c4
+ bl_int_29_4 bl_int_28_4 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c5
+ bl_int_29_5 bl_int_28_5 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c6
+ bl_int_29_6 bl_int_28_6 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c7
+ bl_int_29_7 bl_int_28_7 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c8
+ bl_int_29_8 bl_int_28_8 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c9
+ bl_int_29_9 bl_int_28_9 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c10
+ bl_int_29_10 bl_int_28_10 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c11
+ bl_int_29_11 bl_int_28_11 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c12
+ bl_int_29_12 bl_int_28_12 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c13
+ bl_int_29_13 bl_int_28_13 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c14
+ bl_int_29_14 bl_int_28_14 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c15
+ bl_int_29_15 bl_int_28_15 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c16
+ bl_int_29_16 bl_int_28_16 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c17
+ bl_int_29_17 bl_int_28_17 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c18
+ bl_int_29_18 bl_int_28_18 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c19
+ bl_int_29_19 bl_int_28_19 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c20
+ bl_int_29_20 bl_int_28_20 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c21
+ bl_int_29_21 bl_int_28_21 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c22
+ bl_int_29_22 bl_int_28_22 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c23
+ bl_int_29_23 bl_int_28_23 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c24
+ bl_int_29_24 bl_int_28_24 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c25
+ bl_int_29_25 bl_int_28_25 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c26
+ bl_int_29_26 bl_int_28_26 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c27
+ bl_int_29_27 bl_int_28_27 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c28
+ bl_int_29_28 bl_int_28_28 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c29
+ bl_int_29_29 bl_int_28_29 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c30
+ bl_int_29_30 bl_int_28_30 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c31
+ bl_int_29_31 bl_int_28_31 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c32
+ bl_int_29_32 bl_int_28_32 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c33
+ bl_int_29_33 bl_int_28_33 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c34
+ bl_int_29_34 bl_int_28_34 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c35
+ bl_int_29_35 bl_int_28_35 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c36
+ bl_int_29_36 bl_int_28_36 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c37
+ bl_int_29_37 bl_int_28_37 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c38
+ bl_int_29_38 bl_int_28_38 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c39
+ bl_int_29_39 bl_int_28_39 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c40
+ bl_int_29_40 bl_int_28_40 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c41
+ bl_int_29_41 bl_int_28_41 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c42
+ bl_int_29_42 bl_int_28_42 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c43
+ bl_int_29_43 bl_int_28_43 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c44
+ bl_int_29_44 bl_int_28_44 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c45
+ bl_int_29_45 bl_int_28_45 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c46
+ bl_int_29_46 bl_int_28_46 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c47
+ bl_int_29_47 bl_int_28_47 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c48
+ bl_int_29_48 bl_int_28_48 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c49
+ bl_int_29_49 bl_int_28_49 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c50
+ bl_int_29_50 bl_int_28_50 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c51
+ bl_int_29_51 bl_int_28_51 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c52
+ bl_int_29_52 bl_int_28_52 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c53
+ bl_int_29_53 bl_int_28_53 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c54
+ bl_int_29_54 bl_int_28_54 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c55
+ bl_int_29_55 bl_int_28_55 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c56
+ bl_int_29_56 bl_int_28_56 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c57
+ bl_int_29_57 bl_int_28_57 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c58
+ bl_int_29_58 bl_int_28_58 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c59
+ bl_int_29_59 bl_int_28_59 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c60
+ bl_int_29_60 bl_int_28_60 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c61
+ bl_int_29_61 bl_int_28_61 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c62
+ bl_int_29_62 bl_int_28_62 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c63
+ bl_int_29_63 bl_int_28_63 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c64
+ bl_int_29_64 bl_int_28_64 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c65
+ bl_int_29_65 bl_int_28_65 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c66
+ bl_int_29_66 bl_int_28_66 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c67
+ bl_int_29_67 bl_int_28_67 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c68
+ bl_int_29_68 bl_int_28_68 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c69
+ bl_int_29_69 bl_int_28_69 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c70
+ bl_int_29_70 bl_int_28_70 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c71
+ bl_int_29_71 bl_int_28_71 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c72
+ bl_int_29_72 bl_int_28_72 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c73
+ bl_int_29_73 bl_int_28_73 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c74
+ bl_int_29_74 bl_int_28_74 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c75
+ bl_int_29_75 bl_int_28_75 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c76
+ bl_int_29_76 bl_int_28_76 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c77
+ bl_int_29_77 bl_int_28_77 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c78
+ bl_int_29_78 bl_int_28_78 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c79
+ bl_int_29_79 bl_int_28_79 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c80
+ bl_int_29_80 bl_int_28_80 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c81
+ bl_int_29_81 bl_int_28_81 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c82
+ bl_int_29_82 bl_int_28_82 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c83
+ bl_int_29_83 bl_int_28_83 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c84
+ bl_int_29_84 bl_int_28_84 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c85
+ bl_int_29_85 bl_int_28_85 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c86
+ bl_int_29_86 bl_int_28_86 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c87
+ bl_int_29_87 bl_int_28_87 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c88
+ bl_int_29_88 bl_int_28_88 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c89
+ bl_int_29_89 bl_int_28_89 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c90
+ bl_int_29_90 bl_int_28_90 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c91
+ bl_int_29_91 bl_int_28_91 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c92
+ bl_int_29_92 bl_int_28_92 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c93
+ bl_int_29_93 bl_int_28_93 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c94
+ bl_int_29_94 bl_int_28_94 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c95
+ bl_int_29_95 bl_int_28_95 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c96
+ bl_int_29_96 bl_int_28_96 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c97
+ bl_int_29_97 bl_int_28_97 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c98
+ bl_int_29_98 bl_int_28_98 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c99
+ bl_int_29_99 bl_int_28_99 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c100
+ bl_int_29_100 bl_int_28_100 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c101
+ bl_int_29_101 bl_int_28_101 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c102
+ bl_int_29_102 bl_int_28_102 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c103
+ bl_int_29_103 bl_int_28_103 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c104
+ bl_int_29_104 bl_int_28_104 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c105
+ bl_int_29_105 bl_int_28_105 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c106
+ bl_int_29_106 bl_int_28_106 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c107
+ bl_int_29_107 bl_int_28_107 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c108
+ bl_int_29_108 bl_int_28_108 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c109
+ bl_int_29_109 bl_int_28_109 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c110
+ bl_int_29_110 bl_int_28_110 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c111
+ bl_int_29_111 bl_int_28_111 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c112
+ bl_int_29_112 bl_int_28_112 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c113
+ bl_int_29_113 bl_int_28_113 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c114
+ bl_int_29_114 bl_int_28_114 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c115
+ bl_int_29_115 bl_int_28_115 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c116
+ bl_int_29_116 bl_int_28_116 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c117
+ bl_int_29_117 bl_int_28_117 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c118
+ bl_int_29_118 bl_int_28_118 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c119
+ bl_int_29_119 bl_int_28_119 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c120
+ bl_int_29_120 bl_int_28_120 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c121
+ bl_int_29_121 bl_int_28_121 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c122
+ bl_int_29_122 bl_int_28_122 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c123
+ bl_int_29_123 bl_int_28_123 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c124
+ bl_int_29_124 bl_int_28_124 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c125
+ bl_int_29_125 bl_int_28_125 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c126
+ bl_int_29_126 bl_int_28_126 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c127
+ bl_int_29_127 bl_int_28_127 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c128
+ bl_int_29_128 bl_int_28_128 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c129
+ bl_int_29_129 bl_int_28_129 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c130
+ bl_int_29_130 bl_int_28_130 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c131
+ bl_int_29_131 bl_int_28_131 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c132
+ bl_int_29_132 bl_int_28_132 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c133
+ bl_int_29_133 bl_int_28_133 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c134
+ bl_int_29_134 bl_int_28_134 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c135
+ bl_int_29_135 bl_int_28_135 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c136
+ bl_int_29_136 bl_int_28_136 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c137
+ bl_int_29_137 bl_int_28_137 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c138
+ bl_int_29_138 bl_int_28_138 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c139
+ bl_int_29_139 bl_int_28_139 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c140
+ bl_int_29_140 bl_int_28_140 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c141
+ bl_int_29_141 bl_int_28_141 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c142
+ bl_int_29_142 bl_int_28_142 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c143
+ bl_int_29_143 bl_int_28_143 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c144
+ bl_int_29_144 bl_int_28_144 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c145
+ bl_int_29_145 bl_int_28_145 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c146
+ bl_int_29_146 bl_int_28_146 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c147
+ bl_int_29_147 bl_int_28_147 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c148
+ bl_int_29_148 bl_int_28_148 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c149
+ bl_int_29_149 bl_int_28_149 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c150
+ bl_int_29_150 bl_int_28_150 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c151
+ bl_int_29_151 bl_int_28_151 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c152
+ bl_int_29_152 bl_int_28_152 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c153
+ bl_int_29_153 bl_int_28_153 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c154
+ bl_int_29_154 bl_int_28_154 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c155
+ bl_int_29_155 bl_int_28_155 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c156
+ bl_int_29_156 bl_int_28_156 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c157
+ bl_int_29_157 bl_int_28_157 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c158
+ bl_int_29_158 bl_int_28_158 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c159
+ bl_int_29_159 bl_int_28_159 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c160
+ bl_int_29_160 bl_int_28_160 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c161
+ bl_int_29_161 bl_int_28_161 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c162
+ bl_int_29_162 bl_int_28_162 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c163
+ bl_int_29_163 bl_int_28_163 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c164
+ bl_int_29_164 bl_int_28_164 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c165
+ bl_int_29_165 bl_int_28_165 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c166
+ bl_int_29_166 bl_int_28_166 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c167
+ bl_int_29_167 bl_int_28_167 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c168
+ bl_int_29_168 bl_int_28_168 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c169
+ bl_int_29_169 bl_int_28_169 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c170
+ bl_int_29_170 bl_int_28_170 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c171
+ bl_int_29_171 bl_int_28_171 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c172
+ bl_int_29_172 bl_int_28_172 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c173
+ bl_int_29_173 bl_int_28_173 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c174
+ bl_int_29_174 bl_int_28_174 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c175
+ bl_int_29_175 bl_int_28_175 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c176
+ bl_int_29_176 bl_int_28_176 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c177
+ bl_int_29_177 bl_int_28_177 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c178
+ bl_int_29_178 bl_int_28_178 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c179
+ bl_int_29_179 bl_int_28_179 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c180
+ bl_int_29_180 bl_int_28_180 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c181
+ bl_int_29_181 bl_int_28_181 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c182
+ bl_int_29_182 bl_int_28_182 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r29_c183
+ bl_int_29_183 bl_int_28_183 wl_0_29 gnd
+ sram_rom_base_one_cell
Xbit_r30_c0
+ bl_int_30_0 bl_int_29_0 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c1
+ bl_int_30_1 bl_int_29_1 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c2
+ bl_int_30_2 bl_int_29_2 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c3
+ bl_int_30_3 bl_int_29_3 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c4
+ bl_int_30_4 bl_int_29_4 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c5
+ bl_int_30_5 bl_int_29_5 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c6
+ bl_int_30_6 bl_int_29_6 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c7
+ bl_int_30_7 bl_int_29_7 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c8
+ bl_int_30_8 bl_int_29_8 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c9
+ bl_int_30_9 bl_int_29_9 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c10
+ bl_int_30_10 bl_int_29_10 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c11
+ bl_int_30_11 bl_int_29_11 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c12
+ bl_int_30_12 bl_int_29_12 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c13
+ bl_int_30_13 bl_int_29_13 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c14
+ bl_int_30_14 bl_int_29_14 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c15
+ bl_int_30_15 bl_int_29_15 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c16
+ bl_int_30_16 bl_int_29_16 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c17
+ bl_int_30_17 bl_int_29_17 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c18
+ bl_int_30_18 bl_int_29_18 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c19
+ bl_int_30_19 bl_int_29_19 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c20
+ bl_int_30_20 bl_int_29_20 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c21
+ bl_int_30_21 bl_int_29_21 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c22
+ bl_int_30_22 bl_int_29_22 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c23
+ bl_int_30_23 bl_int_29_23 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c24
+ bl_int_30_24 bl_int_29_24 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c25
+ bl_int_30_25 bl_int_29_25 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c26
+ bl_int_30_26 bl_int_29_26 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c27
+ bl_int_30_27 bl_int_29_27 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c28
+ bl_int_30_28 bl_int_29_28 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c29
+ bl_int_30_29 bl_int_29_29 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c30
+ bl_int_30_30 bl_int_29_30 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c31
+ bl_int_30_31 bl_int_29_31 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c32
+ bl_int_30_32 bl_int_29_32 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c33
+ bl_int_30_33 bl_int_29_33 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c34
+ bl_int_30_34 bl_int_29_34 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c35
+ bl_int_30_35 bl_int_29_35 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c36
+ bl_int_30_36 bl_int_29_36 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c37
+ bl_int_30_37 bl_int_29_37 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c38
+ bl_int_30_38 bl_int_29_38 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c39
+ bl_int_30_39 bl_int_29_39 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c40
+ bl_int_30_40 bl_int_29_40 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c41
+ bl_int_30_41 bl_int_29_41 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c42
+ bl_int_30_42 bl_int_29_42 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c43
+ bl_int_30_43 bl_int_29_43 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c44
+ bl_int_30_44 bl_int_29_44 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c45
+ bl_int_30_45 bl_int_29_45 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c46
+ bl_int_30_46 bl_int_29_46 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c47
+ bl_int_30_47 bl_int_29_47 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c48
+ bl_int_30_48 bl_int_29_48 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c49
+ bl_int_30_49 bl_int_29_49 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c50
+ bl_int_30_50 bl_int_29_50 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c51
+ bl_int_30_51 bl_int_29_51 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c52
+ bl_int_30_52 bl_int_29_52 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c53
+ bl_int_30_53 bl_int_29_53 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c54
+ bl_int_30_54 bl_int_29_54 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c55
+ bl_int_30_55 bl_int_29_55 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c56
+ bl_int_30_56 bl_int_29_56 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c57
+ bl_int_30_57 bl_int_29_57 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c58
+ bl_int_30_58 bl_int_29_58 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c59
+ bl_int_30_59 bl_int_29_59 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c60
+ bl_int_30_60 bl_int_29_60 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c61
+ bl_int_30_61 bl_int_29_61 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c62
+ bl_int_30_62 bl_int_29_62 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c63
+ bl_int_30_63 bl_int_29_63 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c64
+ bl_int_30_64 bl_int_29_64 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c65
+ bl_int_30_65 bl_int_29_65 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c66
+ bl_int_30_66 bl_int_29_66 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c67
+ bl_int_30_67 bl_int_29_67 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c68
+ bl_int_30_68 bl_int_29_68 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c69
+ bl_int_30_69 bl_int_29_69 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c70
+ bl_int_30_70 bl_int_29_70 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c71
+ bl_int_30_71 bl_int_29_71 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c72
+ bl_int_30_72 bl_int_29_72 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c73
+ bl_int_30_73 bl_int_29_73 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c74
+ bl_int_30_74 bl_int_29_74 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c75
+ bl_int_30_75 bl_int_29_75 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c76
+ bl_int_30_76 bl_int_29_76 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c77
+ bl_int_30_77 bl_int_29_77 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c78
+ bl_int_30_78 bl_int_29_78 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c79
+ bl_int_30_79 bl_int_29_79 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c80
+ bl_int_30_80 bl_int_29_80 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c81
+ bl_int_30_81 bl_int_29_81 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c82
+ bl_int_30_82 bl_int_29_82 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c83
+ bl_int_30_83 bl_int_29_83 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c84
+ bl_int_30_84 bl_int_29_84 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c85
+ bl_int_30_85 bl_int_29_85 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c86
+ bl_int_30_86 bl_int_29_86 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c87
+ bl_int_30_87 bl_int_29_87 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c88
+ bl_int_30_88 bl_int_29_88 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c89
+ bl_int_30_89 bl_int_29_89 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c90
+ bl_int_30_90 bl_int_29_90 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c91
+ bl_int_30_91 bl_int_29_91 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c92
+ bl_int_30_92 bl_int_29_92 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c93
+ bl_int_30_93 bl_int_29_93 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c94
+ bl_int_30_94 bl_int_29_94 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c95
+ bl_int_30_95 bl_int_29_95 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c96
+ bl_int_30_96 bl_int_29_96 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c97
+ bl_int_30_97 bl_int_29_97 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c98
+ bl_int_30_98 bl_int_29_98 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c99
+ bl_int_30_99 bl_int_29_99 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c100
+ bl_int_30_100 bl_int_29_100 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c101
+ bl_int_30_101 bl_int_29_101 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c102
+ bl_int_30_102 bl_int_29_102 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c103
+ bl_int_30_103 bl_int_29_103 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c104
+ bl_int_30_104 bl_int_29_104 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c105
+ bl_int_30_105 bl_int_29_105 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c106
+ bl_int_30_106 bl_int_29_106 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c107
+ bl_int_30_107 bl_int_29_107 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c108
+ bl_int_30_108 bl_int_29_108 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c109
+ bl_int_30_109 bl_int_29_109 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c110
+ bl_int_30_110 bl_int_29_110 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c111
+ bl_int_30_111 bl_int_29_111 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c112
+ bl_int_30_112 bl_int_29_112 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c113
+ bl_int_30_113 bl_int_29_113 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c114
+ bl_int_30_114 bl_int_29_114 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c115
+ bl_int_30_115 bl_int_29_115 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c116
+ bl_int_30_116 bl_int_29_116 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c117
+ bl_int_30_117 bl_int_29_117 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c118
+ bl_int_30_118 bl_int_29_118 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c119
+ bl_int_30_119 bl_int_29_119 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c120
+ bl_int_30_120 bl_int_29_120 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c121
+ bl_int_30_121 bl_int_29_121 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c122
+ bl_int_30_122 bl_int_29_122 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c123
+ bl_int_30_123 bl_int_29_123 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c124
+ bl_int_30_124 bl_int_29_124 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c125
+ bl_int_30_125 bl_int_29_125 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c126
+ bl_int_30_126 bl_int_29_126 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c127
+ bl_int_30_127 bl_int_29_127 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c128
+ bl_int_30_128 bl_int_29_128 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c129
+ bl_int_30_129 bl_int_29_129 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c130
+ bl_int_30_130 bl_int_29_130 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c131
+ bl_int_30_131 bl_int_29_131 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c132
+ bl_int_30_132 bl_int_29_132 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c133
+ bl_int_30_133 bl_int_29_133 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c134
+ bl_int_30_134 bl_int_29_134 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c135
+ bl_int_30_135 bl_int_29_135 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c136
+ bl_int_30_136 bl_int_29_136 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c137
+ bl_int_30_137 bl_int_29_137 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c138
+ bl_int_30_138 bl_int_29_138 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c139
+ bl_int_30_139 bl_int_29_139 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c140
+ bl_int_30_140 bl_int_29_140 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c141
+ bl_int_30_141 bl_int_29_141 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c142
+ bl_int_30_142 bl_int_29_142 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c143
+ bl_int_30_143 bl_int_29_143 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c144
+ bl_int_30_144 bl_int_29_144 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c145
+ bl_int_30_145 bl_int_29_145 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c146
+ bl_int_30_146 bl_int_29_146 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c147
+ bl_int_30_147 bl_int_29_147 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c148
+ bl_int_30_148 bl_int_29_148 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c149
+ bl_int_30_149 bl_int_29_149 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c150
+ bl_int_30_150 bl_int_29_150 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c151
+ bl_int_30_151 bl_int_29_151 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c152
+ bl_int_30_152 bl_int_29_152 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c153
+ bl_int_30_153 bl_int_29_153 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c154
+ bl_int_30_154 bl_int_29_154 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c155
+ bl_int_30_155 bl_int_29_155 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c156
+ bl_int_30_156 bl_int_29_156 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c157
+ bl_int_30_157 bl_int_29_157 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c158
+ bl_int_30_158 bl_int_29_158 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c159
+ bl_int_30_159 bl_int_29_159 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c160
+ bl_int_30_160 bl_int_29_160 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c161
+ bl_int_30_161 bl_int_29_161 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c162
+ bl_int_30_162 bl_int_29_162 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c163
+ bl_int_30_163 bl_int_29_163 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c164
+ bl_int_30_164 bl_int_29_164 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c165
+ bl_int_30_165 bl_int_29_165 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c166
+ bl_int_30_166 bl_int_29_166 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c167
+ bl_int_30_167 bl_int_29_167 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c168
+ bl_int_30_168 bl_int_29_168 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c169
+ bl_int_30_169 bl_int_29_169 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c170
+ bl_int_30_170 bl_int_29_170 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c171
+ bl_int_30_171 bl_int_29_171 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c172
+ bl_int_30_172 bl_int_29_172 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c173
+ bl_int_30_173 bl_int_29_173 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c174
+ bl_int_30_174 bl_int_29_174 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c175
+ bl_int_30_175 bl_int_29_175 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c176
+ bl_int_30_176 bl_int_29_176 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c177
+ bl_int_30_177 bl_int_29_177 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c178
+ bl_int_30_178 bl_int_29_178 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c179
+ bl_int_30_179 bl_int_29_179 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c180
+ bl_int_30_180 bl_int_29_180 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c181
+ bl_int_30_181 bl_int_29_181 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c182
+ bl_int_30_182 bl_int_29_182 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r30_c183
+ bl_int_30_183 bl_int_29_183 wl_0_30 gnd
+ sram_rom_base_one_cell
Xbit_r31_c0
+ bl_int_31_0 bl_int_30_0 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c1
+ bl_int_31_1 bl_int_30_1 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c2
+ bl_int_31_2 bl_int_30_2 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c3
+ bl_int_31_3 bl_int_30_3 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c4
+ bl_int_31_4 bl_int_30_4 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c5
+ bl_int_31_5 bl_int_30_5 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c6
+ bl_int_31_6 bl_int_30_6 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c7
+ bl_int_31_7 bl_int_30_7 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c8
+ bl_int_31_8 bl_int_30_8 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c9
+ bl_int_31_9 bl_int_30_9 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c10
+ bl_int_31_10 bl_int_30_10 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c11
+ bl_int_31_11 bl_int_30_11 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c12
+ bl_int_31_12 bl_int_30_12 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c13
+ bl_int_31_13 bl_int_30_13 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c14
+ bl_int_31_14 bl_int_30_14 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c15
+ bl_int_31_15 bl_int_30_15 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c16
+ bl_int_31_16 bl_int_30_16 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c17
+ bl_int_31_17 bl_int_30_17 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c18
+ bl_int_31_18 bl_int_30_18 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c19
+ bl_int_31_19 bl_int_30_19 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c20
+ bl_int_31_20 bl_int_30_20 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c21
+ bl_int_31_21 bl_int_30_21 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c22
+ bl_int_31_22 bl_int_30_22 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c23
+ bl_int_31_23 bl_int_30_23 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c24
+ bl_int_31_24 bl_int_30_24 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c25
+ bl_int_31_25 bl_int_30_25 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c26
+ bl_int_31_26 bl_int_30_26 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c27
+ bl_int_31_27 bl_int_30_27 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c28
+ bl_int_31_28 bl_int_30_28 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c29
+ bl_int_31_29 bl_int_30_29 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c30
+ bl_int_31_30 bl_int_30_30 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c31
+ bl_int_31_31 bl_int_30_31 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c32
+ bl_int_31_32 bl_int_30_32 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c33
+ bl_int_31_33 bl_int_30_33 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c34
+ bl_int_31_34 bl_int_30_34 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c35
+ bl_int_31_35 bl_int_30_35 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c36
+ bl_int_31_36 bl_int_30_36 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c37
+ bl_int_31_37 bl_int_30_37 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c38
+ bl_int_31_38 bl_int_30_38 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c39
+ bl_int_31_39 bl_int_30_39 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c40
+ bl_int_31_40 bl_int_30_40 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c41
+ bl_int_31_41 bl_int_30_41 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c42
+ bl_int_31_42 bl_int_30_42 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c43
+ bl_int_31_43 bl_int_30_43 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c44
+ bl_int_31_44 bl_int_30_44 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c45
+ bl_int_31_45 bl_int_30_45 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c46
+ bl_int_31_46 bl_int_30_46 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c47
+ bl_int_31_47 bl_int_30_47 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c48
+ bl_int_31_48 bl_int_30_48 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c49
+ bl_int_31_49 bl_int_30_49 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c50
+ bl_int_31_50 bl_int_30_50 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c51
+ bl_int_31_51 bl_int_30_51 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c52
+ bl_int_31_52 bl_int_30_52 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c53
+ bl_int_31_53 bl_int_30_53 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c54
+ bl_int_31_54 bl_int_30_54 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c55
+ bl_int_31_55 bl_int_30_55 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c56
+ bl_int_31_56 bl_int_30_56 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c57
+ bl_int_31_57 bl_int_30_57 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c58
+ bl_int_31_58 bl_int_30_58 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c59
+ bl_int_31_59 bl_int_30_59 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c60
+ bl_int_31_60 bl_int_30_60 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c61
+ bl_int_31_61 bl_int_30_61 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c62
+ bl_int_31_62 bl_int_30_62 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c63
+ bl_int_31_63 bl_int_30_63 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c64
+ bl_int_31_64 bl_int_30_64 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c65
+ bl_int_31_65 bl_int_30_65 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c66
+ bl_int_31_66 bl_int_30_66 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c67
+ bl_int_31_67 bl_int_30_67 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c68
+ bl_int_31_68 bl_int_30_68 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c69
+ bl_int_31_69 bl_int_30_69 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c70
+ bl_int_31_70 bl_int_30_70 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c71
+ bl_int_31_71 bl_int_30_71 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c72
+ bl_int_31_72 bl_int_30_72 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c73
+ bl_int_31_73 bl_int_30_73 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c74
+ bl_int_31_74 bl_int_30_74 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c75
+ bl_int_31_75 bl_int_30_75 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c76
+ bl_int_31_76 bl_int_30_76 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c77
+ bl_int_31_77 bl_int_30_77 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c78
+ bl_int_31_78 bl_int_30_78 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c79
+ bl_int_31_79 bl_int_30_79 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c80
+ bl_int_31_80 bl_int_30_80 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c81
+ bl_int_31_81 bl_int_30_81 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c82
+ bl_int_31_82 bl_int_30_82 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c83
+ bl_int_31_83 bl_int_30_83 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c84
+ bl_int_31_84 bl_int_30_84 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c85
+ bl_int_31_85 bl_int_30_85 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c86
+ bl_int_31_86 bl_int_30_86 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c87
+ bl_int_31_87 bl_int_30_87 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c88
+ bl_int_31_88 bl_int_30_88 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c89
+ bl_int_31_89 bl_int_30_89 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c90
+ bl_int_31_90 bl_int_30_90 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c91
+ bl_int_31_91 bl_int_30_91 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c92
+ bl_int_31_92 bl_int_30_92 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c93
+ bl_int_31_93 bl_int_30_93 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c94
+ bl_int_31_94 bl_int_30_94 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c95
+ bl_int_31_95 bl_int_30_95 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c96
+ bl_int_31_96 bl_int_30_96 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c97
+ bl_int_31_97 bl_int_30_97 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c98
+ bl_int_31_98 bl_int_30_98 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c99
+ bl_int_31_99 bl_int_30_99 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c100
+ bl_int_31_100 bl_int_30_100 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c101
+ bl_int_31_101 bl_int_30_101 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c102
+ bl_int_31_102 bl_int_30_102 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c103
+ bl_int_31_103 bl_int_30_103 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c104
+ bl_int_31_104 bl_int_30_104 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c105
+ bl_int_31_105 bl_int_30_105 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c106
+ bl_int_31_106 bl_int_30_106 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c107
+ bl_int_31_107 bl_int_30_107 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c108
+ bl_int_31_108 bl_int_30_108 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c109
+ bl_int_31_109 bl_int_30_109 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c110
+ bl_int_31_110 bl_int_30_110 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c111
+ bl_int_31_111 bl_int_30_111 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c112
+ bl_int_31_112 bl_int_30_112 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c113
+ bl_int_31_113 bl_int_30_113 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c114
+ bl_int_31_114 bl_int_30_114 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c115
+ bl_int_31_115 bl_int_30_115 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c116
+ bl_int_31_116 bl_int_30_116 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c117
+ bl_int_31_117 bl_int_30_117 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c118
+ bl_int_31_118 bl_int_30_118 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c119
+ bl_int_31_119 bl_int_30_119 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c120
+ bl_int_31_120 bl_int_30_120 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c121
+ bl_int_31_121 bl_int_30_121 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c122
+ bl_int_31_122 bl_int_30_122 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c123
+ bl_int_31_123 bl_int_30_123 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c124
+ bl_int_31_124 bl_int_30_124 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c125
+ bl_int_31_125 bl_int_30_125 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c126
+ bl_int_31_126 bl_int_30_126 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c127
+ bl_int_31_127 bl_int_30_127 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c128
+ bl_int_31_128 bl_int_30_128 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c129
+ bl_int_31_129 bl_int_30_129 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c130
+ bl_int_31_130 bl_int_30_130 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c131
+ bl_int_31_131 bl_int_30_131 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c132
+ bl_int_31_132 bl_int_30_132 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c133
+ bl_int_31_133 bl_int_30_133 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c134
+ bl_int_31_134 bl_int_30_134 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c135
+ bl_int_31_135 bl_int_30_135 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c136
+ bl_int_31_136 bl_int_30_136 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c137
+ bl_int_31_137 bl_int_30_137 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c138
+ bl_int_31_138 bl_int_30_138 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c139
+ bl_int_31_139 bl_int_30_139 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c140
+ bl_int_31_140 bl_int_30_140 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c141
+ bl_int_31_141 bl_int_30_141 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c142
+ bl_int_31_142 bl_int_30_142 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c143
+ bl_int_31_143 bl_int_30_143 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c144
+ bl_int_31_144 bl_int_30_144 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c145
+ bl_int_31_145 bl_int_30_145 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c146
+ bl_int_31_146 bl_int_30_146 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c147
+ bl_int_31_147 bl_int_30_147 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c148
+ bl_int_31_148 bl_int_30_148 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c149
+ bl_int_31_149 bl_int_30_149 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c150
+ bl_int_31_150 bl_int_30_150 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c151
+ bl_int_31_151 bl_int_30_151 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c152
+ bl_int_31_152 bl_int_30_152 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c153
+ bl_int_31_153 bl_int_30_153 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c154
+ bl_int_31_154 bl_int_30_154 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c155
+ bl_int_31_155 bl_int_30_155 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c156
+ bl_int_31_156 bl_int_30_156 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c157
+ bl_int_31_157 bl_int_30_157 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c158
+ bl_int_31_158 bl_int_30_158 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c159
+ bl_int_31_159 bl_int_30_159 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c160
+ bl_int_31_160 bl_int_30_160 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c161
+ bl_int_31_161 bl_int_30_161 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c162
+ bl_int_31_162 bl_int_30_162 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c163
+ bl_int_31_163 bl_int_30_163 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c164
+ bl_int_31_164 bl_int_30_164 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c165
+ bl_int_31_165 bl_int_30_165 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c166
+ bl_int_31_166 bl_int_30_166 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c167
+ bl_int_31_167 bl_int_30_167 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c168
+ bl_int_31_168 bl_int_30_168 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c169
+ bl_int_31_169 bl_int_30_169 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c170
+ bl_int_31_170 bl_int_30_170 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c171
+ bl_int_31_171 bl_int_30_171 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c172
+ bl_int_31_172 bl_int_30_172 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c173
+ bl_int_31_173 bl_int_30_173 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c174
+ bl_int_31_174 bl_int_30_174 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c175
+ bl_int_31_175 bl_int_30_175 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c176
+ bl_int_31_176 bl_int_30_176 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c177
+ bl_int_31_177 bl_int_30_177 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c178
+ bl_int_31_178 bl_int_30_178 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c179
+ bl_int_31_179 bl_int_30_179 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c180
+ bl_int_31_180 bl_int_30_180 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c181
+ bl_int_31_181 bl_int_30_181 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c182
+ bl_int_31_182 bl_int_30_182 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r31_c183
+ bl_int_31_183 bl_int_30_183 wl_0_31 gnd
+ sram_rom_base_one_cell
Xbit_r32_c0
+ bl_int_32_0 bl_int_31_0 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c1
+ bl_int_32_1 bl_int_31_1 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c2
+ bl_int_32_2 bl_int_31_2 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c3
+ bl_int_32_3 bl_int_31_3 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c4
+ bl_int_32_4 bl_int_31_4 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c5
+ bl_int_32_5 bl_int_31_5 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c6
+ bl_int_32_6 bl_int_31_6 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c7
+ bl_int_32_7 bl_int_31_7 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c8
+ bl_int_32_8 bl_int_31_8 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c9
+ bl_int_32_9 bl_int_31_9 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c10
+ bl_int_32_10 bl_int_31_10 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c11
+ bl_int_32_11 bl_int_31_11 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c12
+ bl_int_32_12 bl_int_31_12 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c13
+ bl_int_32_13 bl_int_31_13 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c14
+ bl_int_32_14 bl_int_31_14 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c15
+ bl_int_32_15 bl_int_31_15 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c16
+ bl_int_32_16 bl_int_31_16 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c17
+ bl_int_32_17 bl_int_31_17 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c18
+ bl_int_32_18 bl_int_31_18 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c19
+ bl_int_32_19 bl_int_31_19 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c20
+ bl_int_32_20 bl_int_31_20 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c21
+ bl_int_32_21 bl_int_31_21 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c22
+ bl_int_32_22 bl_int_31_22 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c23
+ bl_int_32_23 bl_int_31_23 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c24
+ bl_int_32_24 bl_int_31_24 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c25
+ bl_int_32_25 bl_int_31_25 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c26
+ bl_int_32_26 bl_int_31_26 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c27
+ bl_int_32_27 bl_int_31_27 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c28
+ bl_int_32_28 bl_int_31_28 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c29
+ bl_int_32_29 bl_int_31_29 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c30
+ bl_int_32_30 bl_int_31_30 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c31
+ bl_int_32_31 bl_int_31_31 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c32
+ bl_int_32_32 bl_int_31_32 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c33
+ bl_int_32_33 bl_int_31_33 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c34
+ bl_int_32_34 bl_int_31_34 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c35
+ bl_int_32_35 bl_int_31_35 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c36
+ bl_int_32_36 bl_int_31_36 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c37
+ bl_int_32_37 bl_int_31_37 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c38
+ bl_int_32_38 bl_int_31_38 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c39
+ bl_int_32_39 bl_int_31_39 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c40
+ bl_int_32_40 bl_int_31_40 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c41
+ bl_int_32_41 bl_int_31_41 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c42
+ bl_int_32_42 bl_int_31_42 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c43
+ bl_int_32_43 bl_int_31_43 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c44
+ bl_int_32_44 bl_int_31_44 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c45
+ bl_int_32_45 bl_int_31_45 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c46
+ bl_int_32_46 bl_int_31_46 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c47
+ bl_int_32_47 bl_int_31_47 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c48
+ bl_int_32_48 bl_int_31_48 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c49
+ bl_int_32_49 bl_int_31_49 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c50
+ bl_int_32_50 bl_int_31_50 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c51
+ bl_int_32_51 bl_int_31_51 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c52
+ bl_int_32_52 bl_int_31_52 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c53
+ bl_int_32_53 bl_int_31_53 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c54
+ bl_int_32_54 bl_int_31_54 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c55
+ bl_int_32_55 bl_int_31_55 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c56
+ bl_int_32_56 bl_int_31_56 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c57
+ bl_int_32_57 bl_int_31_57 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c58
+ bl_int_32_58 bl_int_31_58 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c59
+ bl_int_32_59 bl_int_31_59 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c60
+ bl_int_32_60 bl_int_31_60 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c61
+ bl_int_32_61 bl_int_31_61 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c62
+ bl_int_32_62 bl_int_31_62 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c63
+ bl_int_32_63 bl_int_31_63 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c64
+ bl_int_32_64 bl_int_31_64 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c65
+ bl_int_32_65 bl_int_31_65 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c66
+ bl_int_32_66 bl_int_31_66 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c67
+ bl_int_32_67 bl_int_31_67 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c68
+ bl_int_32_68 bl_int_31_68 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c69
+ bl_int_32_69 bl_int_31_69 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c70
+ bl_int_32_70 bl_int_31_70 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c71
+ bl_int_32_71 bl_int_31_71 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c72
+ bl_int_32_72 bl_int_31_72 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c73
+ bl_int_32_73 bl_int_31_73 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c74
+ bl_int_32_74 bl_int_31_74 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c75
+ bl_int_32_75 bl_int_31_75 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c76
+ bl_int_32_76 bl_int_31_76 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c77
+ bl_int_32_77 bl_int_31_77 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c78
+ bl_int_32_78 bl_int_31_78 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c79
+ bl_int_32_79 bl_int_31_79 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c80
+ bl_int_32_80 bl_int_31_80 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c81
+ bl_int_32_81 bl_int_31_81 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c82
+ bl_int_32_82 bl_int_31_82 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c83
+ bl_int_32_83 bl_int_31_83 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c84
+ bl_int_32_84 bl_int_31_84 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c85
+ bl_int_32_85 bl_int_31_85 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c86
+ bl_int_32_86 bl_int_31_86 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c87
+ bl_int_32_87 bl_int_31_87 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c88
+ bl_int_32_88 bl_int_31_88 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c89
+ bl_int_32_89 bl_int_31_89 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c90
+ bl_int_32_90 bl_int_31_90 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c91
+ bl_int_32_91 bl_int_31_91 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c92
+ bl_int_32_92 bl_int_31_92 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c93
+ bl_int_32_93 bl_int_31_93 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c94
+ bl_int_32_94 bl_int_31_94 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c95
+ bl_int_32_95 bl_int_31_95 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c96
+ bl_int_32_96 bl_int_31_96 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c97
+ bl_int_32_97 bl_int_31_97 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c98
+ bl_int_32_98 bl_int_31_98 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c99
+ bl_int_32_99 bl_int_31_99 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c100
+ bl_int_32_100 bl_int_31_100 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c101
+ bl_int_32_101 bl_int_31_101 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c102
+ bl_int_32_102 bl_int_31_102 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c103
+ bl_int_32_103 bl_int_31_103 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c104
+ bl_int_32_104 bl_int_31_104 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c105
+ bl_int_32_105 bl_int_31_105 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c106
+ bl_int_32_106 bl_int_31_106 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c107
+ bl_int_32_107 bl_int_31_107 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c108
+ bl_int_32_108 bl_int_31_108 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c109
+ bl_int_32_109 bl_int_31_109 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c110
+ bl_int_32_110 bl_int_31_110 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c111
+ bl_int_32_111 bl_int_31_111 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c112
+ bl_int_32_112 bl_int_31_112 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c113
+ bl_int_32_113 bl_int_31_113 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c114
+ bl_int_32_114 bl_int_31_114 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c115
+ bl_int_32_115 bl_int_31_115 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c116
+ bl_int_32_116 bl_int_31_116 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c117
+ bl_int_32_117 bl_int_31_117 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c118
+ bl_int_32_118 bl_int_31_118 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c119
+ bl_int_32_119 bl_int_31_119 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c120
+ bl_int_32_120 bl_int_31_120 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c121
+ bl_int_32_121 bl_int_31_121 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c122
+ bl_int_32_122 bl_int_31_122 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c123
+ bl_int_32_123 bl_int_31_123 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c124
+ bl_int_32_124 bl_int_31_124 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c125
+ bl_int_32_125 bl_int_31_125 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c126
+ bl_int_32_126 bl_int_31_126 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c127
+ bl_int_32_127 bl_int_31_127 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c128
+ bl_int_32_128 bl_int_31_128 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c129
+ bl_int_32_129 bl_int_31_129 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c130
+ bl_int_32_130 bl_int_31_130 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c131
+ bl_int_32_131 bl_int_31_131 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c132
+ bl_int_32_132 bl_int_31_132 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c133
+ bl_int_32_133 bl_int_31_133 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c134
+ bl_int_32_134 bl_int_31_134 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c135
+ bl_int_32_135 bl_int_31_135 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c136
+ bl_int_32_136 bl_int_31_136 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c137
+ bl_int_32_137 bl_int_31_137 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c138
+ bl_int_32_138 bl_int_31_138 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c139
+ bl_int_32_139 bl_int_31_139 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c140
+ bl_int_32_140 bl_int_31_140 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c141
+ bl_int_32_141 bl_int_31_141 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c142
+ bl_int_32_142 bl_int_31_142 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c143
+ bl_int_32_143 bl_int_31_143 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c144
+ bl_int_32_144 bl_int_31_144 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c145
+ bl_int_32_145 bl_int_31_145 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c146
+ bl_int_32_146 bl_int_31_146 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c147
+ bl_int_32_147 bl_int_31_147 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c148
+ bl_int_32_148 bl_int_31_148 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c149
+ bl_int_32_149 bl_int_31_149 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c150
+ bl_int_32_150 bl_int_31_150 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c151
+ bl_int_32_151 bl_int_31_151 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c152
+ bl_int_32_152 bl_int_31_152 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c153
+ bl_int_32_153 bl_int_31_153 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c154
+ bl_int_32_154 bl_int_31_154 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c155
+ bl_int_32_155 bl_int_31_155 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c156
+ bl_int_32_156 bl_int_31_156 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c157
+ bl_int_32_157 bl_int_31_157 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c158
+ bl_int_32_158 bl_int_31_158 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c159
+ bl_int_32_159 bl_int_31_159 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c160
+ bl_int_32_160 bl_int_31_160 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c161
+ bl_int_32_161 bl_int_31_161 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c162
+ bl_int_32_162 bl_int_31_162 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c163
+ bl_int_32_163 bl_int_31_163 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c164
+ bl_int_32_164 bl_int_31_164 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c165
+ bl_int_32_165 bl_int_31_165 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c166
+ bl_int_32_166 bl_int_31_166 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c167
+ bl_int_32_167 bl_int_31_167 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c168
+ bl_int_32_168 bl_int_31_168 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c169
+ bl_int_32_169 bl_int_31_169 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c170
+ bl_int_32_170 bl_int_31_170 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c171
+ bl_int_32_171 bl_int_31_171 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c172
+ bl_int_32_172 bl_int_31_172 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c173
+ bl_int_32_173 bl_int_31_173 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c174
+ bl_int_32_174 bl_int_31_174 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c175
+ bl_int_32_175 bl_int_31_175 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c176
+ bl_int_32_176 bl_int_31_176 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c177
+ bl_int_32_177 bl_int_31_177 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c178
+ bl_int_32_178 bl_int_31_178 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c179
+ bl_int_32_179 bl_int_31_179 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c180
+ bl_int_32_180 bl_int_31_180 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c181
+ bl_int_32_181 bl_int_31_181 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c182
+ bl_int_32_182 bl_int_31_182 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r32_c183
+ bl_int_32_183 bl_int_31_183 wl_0_32 gnd
+ sram_rom_base_one_cell
Xbit_r33_c0
+ bl_int_33_0 bl_int_32_0 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c1
+ bl_int_33_1 bl_int_32_1 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c2
+ bl_int_33_2 bl_int_32_2 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c3
+ bl_int_33_3 bl_int_32_3 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c4
+ bl_int_33_4 bl_int_32_4 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c5
+ bl_int_33_5 bl_int_32_5 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c6
+ bl_int_33_6 bl_int_32_6 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c7
+ bl_int_33_7 bl_int_32_7 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c8
+ bl_int_33_8 bl_int_32_8 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c9
+ bl_int_33_9 bl_int_32_9 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c10
+ bl_int_33_10 bl_int_32_10 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c11
+ bl_int_33_11 bl_int_32_11 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c12
+ bl_int_33_12 bl_int_32_12 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c13
+ bl_int_33_13 bl_int_32_13 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c14
+ bl_int_33_14 bl_int_32_14 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c15
+ bl_int_33_15 bl_int_32_15 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c16
+ bl_int_33_16 bl_int_32_16 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c17
+ bl_int_33_17 bl_int_32_17 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c18
+ bl_int_33_18 bl_int_32_18 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c19
+ bl_int_33_19 bl_int_32_19 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c20
+ bl_int_33_20 bl_int_32_20 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c21
+ bl_int_33_21 bl_int_32_21 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c22
+ bl_int_33_22 bl_int_32_22 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c23
+ bl_int_33_23 bl_int_32_23 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c24
+ bl_int_33_24 bl_int_32_24 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c25
+ bl_int_33_25 bl_int_32_25 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c26
+ bl_int_33_26 bl_int_32_26 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c27
+ bl_int_33_27 bl_int_32_27 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c28
+ bl_int_33_28 bl_int_32_28 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c29
+ bl_int_33_29 bl_int_32_29 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c30
+ bl_int_33_30 bl_int_32_30 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c31
+ bl_int_33_31 bl_int_32_31 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c32
+ bl_int_33_32 bl_int_32_32 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c33
+ bl_int_33_33 bl_int_32_33 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c34
+ bl_int_33_34 bl_int_32_34 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c35
+ bl_int_33_35 bl_int_32_35 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c36
+ bl_int_33_36 bl_int_32_36 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c37
+ bl_int_33_37 bl_int_32_37 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c38
+ bl_int_33_38 bl_int_32_38 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c39
+ bl_int_33_39 bl_int_32_39 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c40
+ bl_int_33_40 bl_int_32_40 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c41
+ bl_int_33_41 bl_int_32_41 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c42
+ bl_int_33_42 bl_int_32_42 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c43
+ bl_int_33_43 bl_int_32_43 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c44
+ bl_int_33_44 bl_int_32_44 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c45
+ bl_int_33_45 bl_int_32_45 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c46
+ bl_int_33_46 bl_int_32_46 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c47
+ bl_int_33_47 bl_int_32_47 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c48
+ bl_int_33_48 bl_int_32_48 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c49
+ bl_int_33_49 bl_int_32_49 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c50
+ bl_int_33_50 bl_int_32_50 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c51
+ bl_int_33_51 bl_int_32_51 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c52
+ bl_int_33_52 bl_int_32_52 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c53
+ bl_int_33_53 bl_int_32_53 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c54
+ bl_int_33_54 bl_int_32_54 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c55
+ bl_int_33_55 bl_int_32_55 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c56
+ bl_int_33_56 bl_int_32_56 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c57
+ bl_int_33_57 bl_int_32_57 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c58
+ bl_int_33_58 bl_int_32_58 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c59
+ bl_int_33_59 bl_int_32_59 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c60
+ bl_int_33_60 bl_int_32_60 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c61
+ bl_int_33_61 bl_int_32_61 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c62
+ bl_int_33_62 bl_int_32_62 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c63
+ bl_int_33_63 bl_int_32_63 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c64
+ bl_int_33_64 bl_int_32_64 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c65
+ bl_int_33_65 bl_int_32_65 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c66
+ bl_int_33_66 bl_int_32_66 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c67
+ bl_int_33_67 bl_int_32_67 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c68
+ bl_int_33_68 bl_int_32_68 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c69
+ bl_int_33_69 bl_int_32_69 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c70
+ bl_int_33_70 bl_int_32_70 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c71
+ bl_int_33_71 bl_int_32_71 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c72
+ bl_int_33_72 bl_int_32_72 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c73
+ bl_int_33_73 bl_int_32_73 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c74
+ bl_int_33_74 bl_int_32_74 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c75
+ bl_int_33_75 bl_int_32_75 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c76
+ bl_int_33_76 bl_int_32_76 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c77
+ bl_int_33_77 bl_int_32_77 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c78
+ bl_int_33_78 bl_int_32_78 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c79
+ bl_int_33_79 bl_int_32_79 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c80
+ bl_int_33_80 bl_int_32_80 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c81
+ bl_int_33_81 bl_int_32_81 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c82
+ bl_int_33_82 bl_int_32_82 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c83
+ bl_int_33_83 bl_int_32_83 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c84
+ bl_int_33_84 bl_int_32_84 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c85
+ bl_int_33_85 bl_int_32_85 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c86
+ bl_int_33_86 bl_int_32_86 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c87
+ bl_int_33_87 bl_int_32_87 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c88
+ bl_int_33_88 bl_int_32_88 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c89
+ bl_int_33_89 bl_int_32_89 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c90
+ bl_int_33_90 bl_int_32_90 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c91
+ bl_int_33_91 bl_int_32_91 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c92
+ bl_int_33_92 bl_int_32_92 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c93
+ bl_int_33_93 bl_int_32_93 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c94
+ bl_int_33_94 bl_int_32_94 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c95
+ bl_int_33_95 bl_int_32_95 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c96
+ bl_int_33_96 bl_int_32_96 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c97
+ bl_int_33_97 bl_int_32_97 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c98
+ bl_int_33_98 bl_int_32_98 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c99
+ bl_int_33_99 bl_int_32_99 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c100
+ bl_int_33_100 bl_int_32_100 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c101
+ bl_int_33_101 bl_int_32_101 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c102
+ bl_int_33_102 bl_int_32_102 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c103
+ bl_int_33_103 bl_int_32_103 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c104
+ bl_int_33_104 bl_int_32_104 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c105
+ bl_int_33_105 bl_int_32_105 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c106
+ bl_int_33_106 bl_int_32_106 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c107
+ bl_int_33_107 bl_int_32_107 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c108
+ bl_int_33_108 bl_int_32_108 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c109
+ bl_int_33_109 bl_int_32_109 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c110
+ bl_int_33_110 bl_int_32_110 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c111
+ bl_int_33_111 bl_int_32_111 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c112
+ bl_int_33_112 bl_int_32_112 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c113
+ bl_int_33_113 bl_int_32_113 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c114
+ bl_int_33_114 bl_int_32_114 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c115
+ bl_int_33_115 bl_int_32_115 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c116
+ bl_int_33_116 bl_int_32_116 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c117
+ bl_int_33_117 bl_int_32_117 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c118
+ bl_int_33_118 bl_int_32_118 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c119
+ bl_int_33_119 bl_int_32_119 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c120
+ bl_int_33_120 bl_int_32_120 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c121
+ bl_int_33_121 bl_int_32_121 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c122
+ bl_int_33_122 bl_int_32_122 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c123
+ bl_int_33_123 bl_int_32_123 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c124
+ bl_int_33_124 bl_int_32_124 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c125
+ bl_int_33_125 bl_int_32_125 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c126
+ bl_int_33_126 bl_int_32_126 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c127
+ bl_int_33_127 bl_int_32_127 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c128
+ bl_int_33_128 bl_int_32_128 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c129
+ bl_int_33_129 bl_int_32_129 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c130
+ bl_int_33_130 bl_int_32_130 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c131
+ bl_int_33_131 bl_int_32_131 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c132
+ bl_int_33_132 bl_int_32_132 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c133
+ bl_int_33_133 bl_int_32_133 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c134
+ bl_int_33_134 bl_int_32_134 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c135
+ bl_int_33_135 bl_int_32_135 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c136
+ bl_int_33_136 bl_int_32_136 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c137
+ bl_int_33_137 bl_int_32_137 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c138
+ bl_int_33_138 bl_int_32_138 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c139
+ bl_int_33_139 bl_int_32_139 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c140
+ bl_int_33_140 bl_int_32_140 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c141
+ bl_int_33_141 bl_int_32_141 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c142
+ bl_int_33_142 bl_int_32_142 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c143
+ bl_int_33_143 bl_int_32_143 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c144
+ bl_int_33_144 bl_int_32_144 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c145
+ bl_int_33_145 bl_int_32_145 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c146
+ bl_int_33_146 bl_int_32_146 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c147
+ bl_int_33_147 bl_int_32_147 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c148
+ bl_int_33_148 bl_int_32_148 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c149
+ bl_int_33_149 bl_int_32_149 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c150
+ bl_int_33_150 bl_int_32_150 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c151
+ bl_int_33_151 bl_int_32_151 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c152
+ bl_int_33_152 bl_int_32_152 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c153
+ bl_int_33_153 bl_int_32_153 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c154
+ bl_int_33_154 bl_int_32_154 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c155
+ bl_int_33_155 bl_int_32_155 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c156
+ bl_int_33_156 bl_int_32_156 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c157
+ bl_int_33_157 bl_int_32_157 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c158
+ bl_int_33_158 bl_int_32_158 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c159
+ bl_int_33_159 bl_int_32_159 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c160
+ bl_int_33_160 bl_int_32_160 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c161
+ bl_int_33_161 bl_int_32_161 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c162
+ bl_int_33_162 bl_int_32_162 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c163
+ bl_int_33_163 bl_int_32_163 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c164
+ bl_int_33_164 bl_int_32_164 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c165
+ bl_int_33_165 bl_int_32_165 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c166
+ bl_int_33_166 bl_int_32_166 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c167
+ bl_int_33_167 bl_int_32_167 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c168
+ bl_int_33_168 bl_int_32_168 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c169
+ bl_int_33_169 bl_int_32_169 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c170
+ bl_int_33_170 bl_int_32_170 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c171
+ bl_int_33_171 bl_int_32_171 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c172
+ bl_int_33_172 bl_int_32_172 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c173
+ bl_int_33_173 bl_int_32_173 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c174
+ bl_int_33_174 bl_int_32_174 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c175
+ bl_int_33_175 bl_int_32_175 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c176
+ bl_int_33_176 bl_int_32_176 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c177
+ bl_int_33_177 bl_int_32_177 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c178
+ bl_int_33_178 bl_int_32_178 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c179
+ bl_int_33_179 bl_int_32_179 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c180
+ bl_int_33_180 bl_int_32_180 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c181
+ bl_int_33_181 bl_int_32_181 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c182
+ bl_int_33_182 bl_int_32_182 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r33_c183
+ bl_int_33_183 bl_int_32_183 wl_0_33 gnd
+ sram_rom_base_one_cell
Xbit_r34_c0
+ bl_int_34_0 bl_int_33_0 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c1
+ bl_int_34_1 bl_int_33_1 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c2
+ bl_int_34_2 bl_int_33_2 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c3
+ bl_int_34_3 bl_int_33_3 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c4
+ bl_int_34_4 bl_int_33_4 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c5
+ bl_int_34_5 bl_int_33_5 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c6
+ bl_int_34_6 bl_int_33_6 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c7
+ bl_int_34_7 bl_int_33_7 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c8
+ bl_int_34_8 bl_int_33_8 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c9
+ bl_int_34_9 bl_int_33_9 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c10
+ bl_int_34_10 bl_int_33_10 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c11
+ bl_int_34_11 bl_int_33_11 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c12
+ bl_int_34_12 bl_int_33_12 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c13
+ bl_int_34_13 bl_int_33_13 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c14
+ bl_int_34_14 bl_int_33_14 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c15
+ bl_int_34_15 bl_int_33_15 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c16
+ bl_int_34_16 bl_int_33_16 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c17
+ bl_int_34_17 bl_int_33_17 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c18
+ bl_int_34_18 bl_int_33_18 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c19
+ bl_int_34_19 bl_int_33_19 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c20
+ bl_int_34_20 bl_int_33_20 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c21
+ bl_int_34_21 bl_int_33_21 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c22
+ bl_int_34_22 bl_int_33_22 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c23
+ bl_int_34_23 bl_int_33_23 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c24
+ bl_int_34_24 bl_int_33_24 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c25
+ bl_int_34_25 bl_int_33_25 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c26
+ bl_int_34_26 bl_int_33_26 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c27
+ bl_int_34_27 bl_int_33_27 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c28
+ bl_int_34_28 bl_int_33_28 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c29
+ bl_int_34_29 bl_int_33_29 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c30
+ bl_int_34_30 bl_int_33_30 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c31
+ bl_int_34_31 bl_int_33_31 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c32
+ bl_int_34_32 bl_int_33_32 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c33
+ bl_int_34_33 bl_int_33_33 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c34
+ bl_int_34_34 bl_int_33_34 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c35
+ bl_int_34_35 bl_int_33_35 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c36
+ bl_int_34_36 bl_int_33_36 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c37
+ bl_int_34_37 bl_int_33_37 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c38
+ bl_int_34_38 bl_int_33_38 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c39
+ bl_int_34_39 bl_int_33_39 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c40
+ bl_int_34_40 bl_int_33_40 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c41
+ bl_int_34_41 bl_int_33_41 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c42
+ bl_int_34_42 bl_int_33_42 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c43
+ bl_int_34_43 bl_int_33_43 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c44
+ bl_int_34_44 bl_int_33_44 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c45
+ bl_int_34_45 bl_int_33_45 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c46
+ bl_int_34_46 bl_int_33_46 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c47
+ bl_int_34_47 bl_int_33_47 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c48
+ bl_int_34_48 bl_int_33_48 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c49
+ bl_int_34_49 bl_int_33_49 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c50
+ bl_int_34_50 bl_int_33_50 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c51
+ bl_int_34_51 bl_int_33_51 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c52
+ bl_int_34_52 bl_int_33_52 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c53
+ bl_int_34_53 bl_int_33_53 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c54
+ bl_int_34_54 bl_int_33_54 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c55
+ bl_int_34_55 bl_int_33_55 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c56
+ bl_int_34_56 bl_int_33_56 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c57
+ bl_int_34_57 bl_int_33_57 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c58
+ bl_int_34_58 bl_int_33_58 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c59
+ bl_int_34_59 bl_int_33_59 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c60
+ bl_int_34_60 bl_int_33_60 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c61
+ bl_int_34_61 bl_int_33_61 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c62
+ bl_int_34_62 bl_int_33_62 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c63
+ bl_int_34_63 bl_int_33_63 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c64
+ bl_int_34_64 bl_int_33_64 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c65
+ bl_int_34_65 bl_int_33_65 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c66
+ bl_int_34_66 bl_int_33_66 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c67
+ bl_int_34_67 bl_int_33_67 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c68
+ bl_int_34_68 bl_int_33_68 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c69
+ bl_int_34_69 bl_int_33_69 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c70
+ bl_int_34_70 bl_int_33_70 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c71
+ bl_int_34_71 bl_int_33_71 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c72
+ bl_int_34_72 bl_int_33_72 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c73
+ bl_int_34_73 bl_int_33_73 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c74
+ bl_int_34_74 bl_int_33_74 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c75
+ bl_int_34_75 bl_int_33_75 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c76
+ bl_int_34_76 bl_int_33_76 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c77
+ bl_int_34_77 bl_int_33_77 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c78
+ bl_int_34_78 bl_int_33_78 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c79
+ bl_int_34_79 bl_int_33_79 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c80
+ bl_int_34_80 bl_int_33_80 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c81
+ bl_int_34_81 bl_int_33_81 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c82
+ bl_int_34_82 bl_int_33_82 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c83
+ bl_int_34_83 bl_int_33_83 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c84
+ bl_int_34_84 bl_int_33_84 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c85
+ bl_int_34_85 bl_int_33_85 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c86
+ bl_int_34_86 bl_int_33_86 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c87
+ bl_int_34_87 bl_int_33_87 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c88
+ bl_int_34_88 bl_int_33_88 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c89
+ bl_int_34_89 bl_int_33_89 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c90
+ bl_int_34_90 bl_int_33_90 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c91
+ bl_int_34_91 bl_int_33_91 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c92
+ bl_int_34_92 bl_int_33_92 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c93
+ bl_int_34_93 bl_int_33_93 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c94
+ bl_int_34_94 bl_int_33_94 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c95
+ bl_int_34_95 bl_int_33_95 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c96
+ bl_int_34_96 bl_int_33_96 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c97
+ bl_int_34_97 bl_int_33_97 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c98
+ bl_int_34_98 bl_int_33_98 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c99
+ bl_int_34_99 bl_int_33_99 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c100
+ bl_int_34_100 bl_int_33_100 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c101
+ bl_int_34_101 bl_int_33_101 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c102
+ bl_int_34_102 bl_int_33_102 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c103
+ bl_int_34_103 bl_int_33_103 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c104
+ bl_int_34_104 bl_int_33_104 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c105
+ bl_int_34_105 bl_int_33_105 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c106
+ bl_int_34_106 bl_int_33_106 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c107
+ bl_int_34_107 bl_int_33_107 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c108
+ bl_int_34_108 bl_int_33_108 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c109
+ bl_int_34_109 bl_int_33_109 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c110
+ bl_int_34_110 bl_int_33_110 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c111
+ bl_int_34_111 bl_int_33_111 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c112
+ bl_int_34_112 bl_int_33_112 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c113
+ bl_int_34_113 bl_int_33_113 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c114
+ bl_int_34_114 bl_int_33_114 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c115
+ bl_int_34_115 bl_int_33_115 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c116
+ bl_int_34_116 bl_int_33_116 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c117
+ bl_int_34_117 bl_int_33_117 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c118
+ bl_int_34_118 bl_int_33_118 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c119
+ bl_int_34_119 bl_int_33_119 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c120
+ bl_int_34_120 bl_int_33_120 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c121
+ bl_int_34_121 bl_int_33_121 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c122
+ bl_int_34_122 bl_int_33_122 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c123
+ bl_int_34_123 bl_int_33_123 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c124
+ bl_int_34_124 bl_int_33_124 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c125
+ bl_int_34_125 bl_int_33_125 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c126
+ bl_int_34_126 bl_int_33_126 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c127
+ bl_int_34_127 bl_int_33_127 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c128
+ bl_int_34_128 bl_int_33_128 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c129
+ bl_int_34_129 bl_int_33_129 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c130
+ bl_int_34_130 bl_int_33_130 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c131
+ bl_int_34_131 bl_int_33_131 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c132
+ bl_int_34_132 bl_int_33_132 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c133
+ bl_int_34_133 bl_int_33_133 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c134
+ bl_int_34_134 bl_int_33_134 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c135
+ bl_int_34_135 bl_int_33_135 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c136
+ bl_int_34_136 bl_int_33_136 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c137
+ bl_int_34_137 bl_int_33_137 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c138
+ bl_int_34_138 bl_int_33_138 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c139
+ bl_int_34_139 bl_int_33_139 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c140
+ bl_int_34_140 bl_int_33_140 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c141
+ bl_int_34_141 bl_int_33_141 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c142
+ bl_int_34_142 bl_int_33_142 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c143
+ bl_int_34_143 bl_int_33_143 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c144
+ bl_int_34_144 bl_int_33_144 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c145
+ bl_int_34_145 bl_int_33_145 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c146
+ bl_int_34_146 bl_int_33_146 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c147
+ bl_int_34_147 bl_int_33_147 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c148
+ bl_int_34_148 bl_int_33_148 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c149
+ bl_int_34_149 bl_int_33_149 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c150
+ bl_int_34_150 bl_int_33_150 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c151
+ bl_int_34_151 bl_int_33_151 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c152
+ bl_int_34_152 bl_int_33_152 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c153
+ bl_int_34_153 bl_int_33_153 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c154
+ bl_int_34_154 bl_int_33_154 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c155
+ bl_int_34_155 bl_int_33_155 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c156
+ bl_int_34_156 bl_int_33_156 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c157
+ bl_int_34_157 bl_int_33_157 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c158
+ bl_int_34_158 bl_int_33_158 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c159
+ bl_int_34_159 bl_int_33_159 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c160
+ bl_int_34_160 bl_int_33_160 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c161
+ bl_int_34_161 bl_int_33_161 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c162
+ bl_int_34_162 bl_int_33_162 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c163
+ bl_int_34_163 bl_int_33_163 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c164
+ bl_int_34_164 bl_int_33_164 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c165
+ bl_int_34_165 bl_int_33_165 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c166
+ bl_int_34_166 bl_int_33_166 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c167
+ bl_int_34_167 bl_int_33_167 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c168
+ bl_int_34_168 bl_int_33_168 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c169
+ bl_int_34_169 bl_int_33_169 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c170
+ bl_int_34_170 bl_int_33_170 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c171
+ bl_int_34_171 bl_int_33_171 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c172
+ bl_int_34_172 bl_int_33_172 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c173
+ bl_int_34_173 bl_int_33_173 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c174
+ bl_int_34_174 bl_int_33_174 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c175
+ bl_int_34_175 bl_int_33_175 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c176
+ bl_int_34_176 bl_int_33_176 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c177
+ bl_int_34_177 bl_int_33_177 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c178
+ bl_int_34_178 bl_int_33_178 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c179
+ bl_int_34_179 bl_int_33_179 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c180
+ bl_int_34_180 bl_int_33_180 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c181
+ bl_int_34_181 bl_int_33_181 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c182
+ bl_int_34_182 bl_int_33_182 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r34_c183
+ bl_int_34_183 bl_int_33_183 wl_0_34 gnd
+ sram_rom_base_one_cell
Xbit_r35_c0
+ bl_int_35_0 bl_int_34_0 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c1
+ bl_int_35_1 bl_int_34_1 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c2
+ bl_int_35_2 bl_int_34_2 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c3
+ bl_int_35_3 bl_int_34_3 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c4
+ bl_int_35_4 bl_int_34_4 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c5
+ bl_int_35_5 bl_int_34_5 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c6
+ bl_int_35_6 bl_int_34_6 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c7
+ bl_int_35_7 bl_int_34_7 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c8
+ bl_int_35_8 bl_int_34_8 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c9
+ bl_int_35_9 bl_int_34_9 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c10
+ bl_int_35_10 bl_int_34_10 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c11
+ bl_int_35_11 bl_int_34_11 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c12
+ bl_int_35_12 bl_int_34_12 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c13
+ bl_int_35_13 bl_int_34_13 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c14
+ bl_int_35_14 bl_int_34_14 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c15
+ bl_int_35_15 bl_int_34_15 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c16
+ bl_int_35_16 bl_int_34_16 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c17
+ bl_int_35_17 bl_int_34_17 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c18
+ bl_int_35_18 bl_int_34_18 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c19
+ bl_int_35_19 bl_int_34_19 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c20
+ bl_int_35_20 bl_int_34_20 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c21
+ bl_int_35_21 bl_int_34_21 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c22
+ bl_int_35_22 bl_int_34_22 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c23
+ bl_int_35_23 bl_int_34_23 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c24
+ bl_int_35_24 bl_int_34_24 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c25
+ bl_int_35_25 bl_int_34_25 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c26
+ bl_int_35_26 bl_int_34_26 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c27
+ bl_int_35_27 bl_int_34_27 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c28
+ bl_int_35_28 bl_int_34_28 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c29
+ bl_int_35_29 bl_int_34_29 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c30
+ bl_int_35_30 bl_int_34_30 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c31
+ bl_int_35_31 bl_int_34_31 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c32
+ bl_int_35_32 bl_int_34_32 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c33
+ bl_int_35_33 bl_int_34_33 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c34
+ bl_int_35_34 bl_int_34_34 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c35
+ bl_int_35_35 bl_int_34_35 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c36
+ bl_int_35_36 bl_int_34_36 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c37
+ bl_int_35_37 bl_int_34_37 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c38
+ bl_int_35_38 bl_int_34_38 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c39
+ bl_int_35_39 bl_int_34_39 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c40
+ bl_int_35_40 bl_int_34_40 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c41
+ bl_int_35_41 bl_int_34_41 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c42
+ bl_int_35_42 bl_int_34_42 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c43
+ bl_int_35_43 bl_int_34_43 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c44
+ bl_int_35_44 bl_int_34_44 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c45
+ bl_int_35_45 bl_int_34_45 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c46
+ bl_int_35_46 bl_int_34_46 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c47
+ bl_int_35_47 bl_int_34_47 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c48
+ bl_int_35_48 bl_int_34_48 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c49
+ bl_int_35_49 bl_int_34_49 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c50
+ bl_int_35_50 bl_int_34_50 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c51
+ bl_int_35_51 bl_int_34_51 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c52
+ bl_int_35_52 bl_int_34_52 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c53
+ bl_int_35_53 bl_int_34_53 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c54
+ bl_int_35_54 bl_int_34_54 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c55
+ bl_int_35_55 bl_int_34_55 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c56
+ bl_int_35_56 bl_int_34_56 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c57
+ bl_int_35_57 bl_int_34_57 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c58
+ bl_int_35_58 bl_int_34_58 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c59
+ bl_int_35_59 bl_int_34_59 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c60
+ bl_int_35_60 bl_int_34_60 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c61
+ bl_int_35_61 bl_int_34_61 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c62
+ bl_int_35_62 bl_int_34_62 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c63
+ bl_int_35_63 bl_int_34_63 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c64
+ bl_int_35_64 bl_int_34_64 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c65
+ bl_int_35_65 bl_int_34_65 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c66
+ bl_int_35_66 bl_int_34_66 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c67
+ bl_int_35_67 bl_int_34_67 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c68
+ bl_int_35_68 bl_int_34_68 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c69
+ bl_int_35_69 bl_int_34_69 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c70
+ bl_int_35_70 bl_int_34_70 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c71
+ bl_int_35_71 bl_int_34_71 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c72
+ bl_int_35_72 bl_int_34_72 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c73
+ bl_int_35_73 bl_int_34_73 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c74
+ bl_int_35_74 bl_int_34_74 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c75
+ bl_int_35_75 bl_int_34_75 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c76
+ bl_int_35_76 bl_int_34_76 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c77
+ bl_int_35_77 bl_int_34_77 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c78
+ bl_int_35_78 bl_int_34_78 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c79
+ bl_int_35_79 bl_int_34_79 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c80
+ bl_int_35_80 bl_int_34_80 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c81
+ bl_int_35_81 bl_int_34_81 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c82
+ bl_int_35_82 bl_int_34_82 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c83
+ bl_int_35_83 bl_int_34_83 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c84
+ bl_int_35_84 bl_int_34_84 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c85
+ bl_int_35_85 bl_int_34_85 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c86
+ bl_int_35_86 bl_int_34_86 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c87
+ bl_int_35_87 bl_int_34_87 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c88
+ bl_int_35_88 bl_int_34_88 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c89
+ bl_int_35_89 bl_int_34_89 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c90
+ bl_int_35_90 bl_int_34_90 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c91
+ bl_int_35_91 bl_int_34_91 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c92
+ bl_int_35_92 bl_int_34_92 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c93
+ bl_int_35_93 bl_int_34_93 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c94
+ bl_int_35_94 bl_int_34_94 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c95
+ bl_int_35_95 bl_int_34_95 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c96
+ bl_int_35_96 bl_int_34_96 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c97
+ bl_int_35_97 bl_int_34_97 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c98
+ bl_int_35_98 bl_int_34_98 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c99
+ bl_int_35_99 bl_int_34_99 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c100
+ bl_int_35_100 bl_int_34_100 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c101
+ bl_int_35_101 bl_int_34_101 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c102
+ bl_int_35_102 bl_int_34_102 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c103
+ bl_int_35_103 bl_int_34_103 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c104
+ bl_int_35_104 bl_int_34_104 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c105
+ bl_int_35_105 bl_int_34_105 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c106
+ bl_int_35_106 bl_int_34_106 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c107
+ bl_int_35_107 bl_int_34_107 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c108
+ bl_int_35_108 bl_int_34_108 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c109
+ bl_int_35_109 bl_int_34_109 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c110
+ bl_int_35_110 bl_int_34_110 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c111
+ bl_int_35_111 bl_int_34_111 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c112
+ bl_int_35_112 bl_int_34_112 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c113
+ bl_int_35_113 bl_int_34_113 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c114
+ bl_int_35_114 bl_int_34_114 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c115
+ bl_int_35_115 bl_int_34_115 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c116
+ bl_int_35_116 bl_int_34_116 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c117
+ bl_int_35_117 bl_int_34_117 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c118
+ bl_int_35_118 bl_int_34_118 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c119
+ bl_int_35_119 bl_int_34_119 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c120
+ bl_int_35_120 bl_int_34_120 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c121
+ bl_int_35_121 bl_int_34_121 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c122
+ bl_int_35_122 bl_int_34_122 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c123
+ bl_int_35_123 bl_int_34_123 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c124
+ bl_int_35_124 bl_int_34_124 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c125
+ bl_int_35_125 bl_int_34_125 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c126
+ bl_int_35_126 bl_int_34_126 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c127
+ bl_int_35_127 bl_int_34_127 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c128
+ bl_int_35_128 bl_int_34_128 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c129
+ bl_int_35_129 bl_int_34_129 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c130
+ bl_int_35_130 bl_int_34_130 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c131
+ bl_int_35_131 bl_int_34_131 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c132
+ bl_int_35_132 bl_int_34_132 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c133
+ bl_int_35_133 bl_int_34_133 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c134
+ bl_int_35_134 bl_int_34_134 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c135
+ bl_int_35_135 bl_int_34_135 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c136
+ bl_int_35_136 bl_int_34_136 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c137
+ bl_int_35_137 bl_int_34_137 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c138
+ bl_int_35_138 bl_int_34_138 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c139
+ bl_int_35_139 bl_int_34_139 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c140
+ bl_int_35_140 bl_int_34_140 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c141
+ bl_int_35_141 bl_int_34_141 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c142
+ bl_int_35_142 bl_int_34_142 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c143
+ bl_int_35_143 bl_int_34_143 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c144
+ bl_int_35_144 bl_int_34_144 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c145
+ bl_int_35_145 bl_int_34_145 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c146
+ bl_int_35_146 bl_int_34_146 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c147
+ bl_int_35_147 bl_int_34_147 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c148
+ bl_int_35_148 bl_int_34_148 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c149
+ bl_int_35_149 bl_int_34_149 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c150
+ bl_int_35_150 bl_int_34_150 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c151
+ bl_int_35_151 bl_int_34_151 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c152
+ bl_int_35_152 bl_int_34_152 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c153
+ bl_int_35_153 bl_int_34_153 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c154
+ bl_int_35_154 bl_int_34_154 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c155
+ bl_int_35_155 bl_int_34_155 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c156
+ bl_int_35_156 bl_int_34_156 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c157
+ bl_int_35_157 bl_int_34_157 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c158
+ bl_int_35_158 bl_int_34_158 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c159
+ bl_int_35_159 bl_int_34_159 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c160
+ bl_int_35_160 bl_int_34_160 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c161
+ bl_int_35_161 bl_int_34_161 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c162
+ bl_int_35_162 bl_int_34_162 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c163
+ bl_int_35_163 bl_int_34_163 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c164
+ bl_int_35_164 bl_int_34_164 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c165
+ bl_int_35_165 bl_int_34_165 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c166
+ bl_int_35_166 bl_int_34_166 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c167
+ bl_int_35_167 bl_int_34_167 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c168
+ bl_int_35_168 bl_int_34_168 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c169
+ bl_int_35_169 bl_int_34_169 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c170
+ bl_int_35_170 bl_int_34_170 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c171
+ bl_int_35_171 bl_int_34_171 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c172
+ bl_int_35_172 bl_int_34_172 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c173
+ bl_int_35_173 bl_int_34_173 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c174
+ bl_int_35_174 bl_int_34_174 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c175
+ bl_int_35_175 bl_int_34_175 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c176
+ bl_int_35_176 bl_int_34_176 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c177
+ bl_int_35_177 bl_int_34_177 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c178
+ bl_int_35_178 bl_int_34_178 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c179
+ bl_int_35_179 bl_int_34_179 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c180
+ bl_int_35_180 bl_int_34_180 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c181
+ bl_int_35_181 bl_int_34_181 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c182
+ bl_int_35_182 bl_int_34_182 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r35_c183
+ bl_int_35_183 bl_int_34_183 wl_0_35 gnd
+ sram_rom_base_one_cell
Xbit_r36_c0
+ bl_int_36_0 bl_int_35_0 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c1
+ bl_int_36_1 bl_int_35_1 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c2
+ bl_int_36_2 bl_int_35_2 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c3
+ bl_int_36_3 bl_int_35_3 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c4
+ bl_int_36_4 bl_int_35_4 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c5
+ bl_int_36_5 bl_int_35_5 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c6
+ bl_int_36_6 bl_int_35_6 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c7
+ bl_int_36_7 bl_int_35_7 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c8
+ bl_int_36_8 bl_int_35_8 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c9
+ bl_int_36_9 bl_int_35_9 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c10
+ bl_int_36_10 bl_int_35_10 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c11
+ bl_int_36_11 bl_int_35_11 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c12
+ bl_int_36_12 bl_int_35_12 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c13
+ bl_int_36_13 bl_int_35_13 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c14
+ bl_int_36_14 bl_int_35_14 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c15
+ bl_int_36_15 bl_int_35_15 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c16
+ bl_int_36_16 bl_int_35_16 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c17
+ bl_int_36_17 bl_int_35_17 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c18
+ bl_int_36_18 bl_int_35_18 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c19
+ bl_int_36_19 bl_int_35_19 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c20
+ bl_int_36_20 bl_int_35_20 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c21
+ bl_int_36_21 bl_int_35_21 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c22
+ bl_int_36_22 bl_int_35_22 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c23
+ bl_int_36_23 bl_int_35_23 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c24
+ bl_int_36_24 bl_int_35_24 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c25
+ bl_int_36_25 bl_int_35_25 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c26
+ bl_int_36_26 bl_int_35_26 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c27
+ bl_int_36_27 bl_int_35_27 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c28
+ bl_int_36_28 bl_int_35_28 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c29
+ bl_int_36_29 bl_int_35_29 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c30
+ bl_int_36_30 bl_int_35_30 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c31
+ bl_int_36_31 bl_int_35_31 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c32
+ bl_int_36_32 bl_int_35_32 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c33
+ bl_int_36_33 bl_int_35_33 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c34
+ bl_int_36_34 bl_int_35_34 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c35
+ bl_int_36_35 bl_int_35_35 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c36
+ bl_int_36_36 bl_int_35_36 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c37
+ bl_int_36_37 bl_int_35_37 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c38
+ bl_int_36_38 bl_int_35_38 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c39
+ bl_int_36_39 bl_int_35_39 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c40
+ bl_int_36_40 bl_int_35_40 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c41
+ bl_int_36_41 bl_int_35_41 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c42
+ bl_int_36_42 bl_int_35_42 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c43
+ bl_int_36_43 bl_int_35_43 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c44
+ bl_int_36_44 bl_int_35_44 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c45
+ bl_int_36_45 bl_int_35_45 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c46
+ bl_int_36_46 bl_int_35_46 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c47
+ bl_int_36_47 bl_int_35_47 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c48
+ bl_int_36_48 bl_int_35_48 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c49
+ bl_int_36_49 bl_int_35_49 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c50
+ bl_int_36_50 bl_int_35_50 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c51
+ bl_int_36_51 bl_int_35_51 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c52
+ bl_int_36_52 bl_int_35_52 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c53
+ bl_int_36_53 bl_int_35_53 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c54
+ bl_int_36_54 bl_int_35_54 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c55
+ bl_int_36_55 bl_int_35_55 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c56
+ bl_int_36_56 bl_int_35_56 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c57
+ bl_int_36_57 bl_int_35_57 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c58
+ bl_int_36_58 bl_int_35_58 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c59
+ bl_int_36_59 bl_int_35_59 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c60
+ bl_int_36_60 bl_int_35_60 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c61
+ bl_int_36_61 bl_int_35_61 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c62
+ bl_int_36_62 bl_int_35_62 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c63
+ bl_int_36_63 bl_int_35_63 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c64
+ bl_int_36_64 bl_int_35_64 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c65
+ bl_int_36_65 bl_int_35_65 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c66
+ bl_int_36_66 bl_int_35_66 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c67
+ bl_int_36_67 bl_int_35_67 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c68
+ bl_int_36_68 bl_int_35_68 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c69
+ bl_int_36_69 bl_int_35_69 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c70
+ bl_int_36_70 bl_int_35_70 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c71
+ bl_int_36_71 bl_int_35_71 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c72
+ bl_int_36_72 bl_int_35_72 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c73
+ bl_int_36_73 bl_int_35_73 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c74
+ bl_int_36_74 bl_int_35_74 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c75
+ bl_int_36_75 bl_int_35_75 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c76
+ bl_int_36_76 bl_int_35_76 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c77
+ bl_int_36_77 bl_int_35_77 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c78
+ bl_int_36_78 bl_int_35_78 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c79
+ bl_int_36_79 bl_int_35_79 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c80
+ bl_int_36_80 bl_int_35_80 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c81
+ bl_int_36_81 bl_int_35_81 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c82
+ bl_int_36_82 bl_int_35_82 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c83
+ bl_int_36_83 bl_int_35_83 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c84
+ bl_int_36_84 bl_int_35_84 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c85
+ bl_int_36_85 bl_int_35_85 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c86
+ bl_int_36_86 bl_int_35_86 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c87
+ bl_int_36_87 bl_int_35_87 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c88
+ bl_int_36_88 bl_int_35_88 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c89
+ bl_int_36_89 bl_int_35_89 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c90
+ bl_int_36_90 bl_int_35_90 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c91
+ bl_int_36_91 bl_int_35_91 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c92
+ bl_int_36_92 bl_int_35_92 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c93
+ bl_int_36_93 bl_int_35_93 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c94
+ bl_int_36_94 bl_int_35_94 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c95
+ bl_int_36_95 bl_int_35_95 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c96
+ bl_int_36_96 bl_int_35_96 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c97
+ bl_int_36_97 bl_int_35_97 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c98
+ bl_int_36_98 bl_int_35_98 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c99
+ bl_int_36_99 bl_int_35_99 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c100
+ bl_int_36_100 bl_int_35_100 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c101
+ bl_int_36_101 bl_int_35_101 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c102
+ bl_int_36_102 bl_int_35_102 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c103
+ bl_int_36_103 bl_int_35_103 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c104
+ bl_int_36_104 bl_int_35_104 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c105
+ bl_int_36_105 bl_int_35_105 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c106
+ bl_int_36_106 bl_int_35_106 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c107
+ bl_int_36_107 bl_int_35_107 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c108
+ bl_int_36_108 bl_int_35_108 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c109
+ bl_int_36_109 bl_int_35_109 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c110
+ bl_int_36_110 bl_int_35_110 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c111
+ bl_int_36_111 bl_int_35_111 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c112
+ bl_int_36_112 bl_int_35_112 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c113
+ bl_int_36_113 bl_int_35_113 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c114
+ bl_int_36_114 bl_int_35_114 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c115
+ bl_int_36_115 bl_int_35_115 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c116
+ bl_int_36_116 bl_int_35_116 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c117
+ bl_int_36_117 bl_int_35_117 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c118
+ bl_int_36_118 bl_int_35_118 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c119
+ bl_int_36_119 bl_int_35_119 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c120
+ bl_int_36_120 bl_int_35_120 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c121
+ bl_int_36_121 bl_int_35_121 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c122
+ bl_int_36_122 bl_int_35_122 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c123
+ bl_int_36_123 bl_int_35_123 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c124
+ bl_int_36_124 bl_int_35_124 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c125
+ bl_int_36_125 bl_int_35_125 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c126
+ bl_int_36_126 bl_int_35_126 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c127
+ bl_int_36_127 bl_int_35_127 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c128
+ bl_int_36_128 bl_int_35_128 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c129
+ bl_int_36_129 bl_int_35_129 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c130
+ bl_int_36_130 bl_int_35_130 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c131
+ bl_int_36_131 bl_int_35_131 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c132
+ bl_int_36_132 bl_int_35_132 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c133
+ bl_int_36_133 bl_int_35_133 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c134
+ bl_int_36_134 bl_int_35_134 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c135
+ bl_int_36_135 bl_int_35_135 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c136
+ bl_int_36_136 bl_int_35_136 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c137
+ bl_int_36_137 bl_int_35_137 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c138
+ bl_int_36_138 bl_int_35_138 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c139
+ bl_int_36_139 bl_int_35_139 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c140
+ bl_int_36_140 bl_int_35_140 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c141
+ bl_int_36_141 bl_int_35_141 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c142
+ bl_int_36_142 bl_int_35_142 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c143
+ bl_int_36_143 bl_int_35_143 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c144
+ bl_int_36_144 bl_int_35_144 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c145
+ bl_int_36_145 bl_int_35_145 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c146
+ bl_int_36_146 bl_int_35_146 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c147
+ bl_int_36_147 bl_int_35_147 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c148
+ bl_int_36_148 bl_int_35_148 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c149
+ bl_int_36_149 bl_int_35_149 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c150
+ bl_int_36_150 bl_int_35_150 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c151
+ bl_int_36_151 bl_int_35_151 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c152
+ bl_int_36_152 bl_int_35_152 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c153
+ bl_int_36_153 bl_int_35_153 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c154
+ bl_int_36_154 bl_int_35_154 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c155
+ bl_int_36_155 bl_int_35_155 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c156
+ bl_int_36_156 bl_int_35_156 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c157
+ bl_int_36_157 bl_int_35_157 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c158
+ bl_int_36_158 bl_int_35_158 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c159
+ bl_int_36_159 bl_int_35_159 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c160
+ bl_int_36_160 bl_int_35_160 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c161
+ bl_int_36_161 bl_int_35_161 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c162
+ bl_int_36_162 bl_int_35_162 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c163
+ bl_int_36_163 bl_int_35_163 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c164
+ bl_int_36_164 bl_int_35_164 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c165
+ bl_int_36_165 bl_int_35_165 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c166
+ bl_int_36_166 bl_int_35_166 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c167
+ bl_int_36_167 bl_int_35_167 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c168
+ bl_int_36_168 bl_int_35_168 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c169
+ bl_int_36_169 bl_int_35_169 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c170
+ bl_int_36_170 bl_int_35_170 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c171
+ bl_int_36_171 bl_int_35_171 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c172
+ bl_int_36_172 bl_int_35_172 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c173
+ bl_int_36_173 bl_int_35_173 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c174
+ bl_int_36_174 bl_int_35_174 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c175
+ bl_int_36_175 bl_int_35_175 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c176
+ bl_int_36_176 bl_int_35_176 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c177
+ bl_int_36_177 bl_int_35_177 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c178
+ bl_int_36_178 bl_int_35_178 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c179
+ bl_int_36_179 bl_int_35_179 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c180
+ bl_int_36_180 bl_int_35_180 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c181
+ bl_int_36_181 bl_int_35_181 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c182
+ bl_int_36_182 bl_int_35_182 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r36_c183
+ bl_int_36_183 bl_int_35_183 wl_0_36 gnd
+ sram_rom_base_one_cell
Xbit_r37_c0
+ bl_int_37_0 bl_int_36_0 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c1
+ bl_int_37_1 bl_int_36_1 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c2
+ bl_int_37_2 bl_int_36_2 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c3
+ bl_int_37_3 bl_int_36_3 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c4
+ bl_int_37_4 bl_int_36_4 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c5
+ bl_int_37_5 bl_int_36_5 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c6
+ bl_int_37_6 bl_int_36_6 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c7
+ bl_int_37_7 bl_int_36_7 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c8
+ bl_int_37_8 bl_int_36_8 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c9
+ bl_int_37_9 bl_int_36_9 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c10
+ bl_int_37_10 bl_int_36_10 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c11
+ bl_int_37_11 bl_int_36_11 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c12
+ bl_int_37_12 bl_int_36_12 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c13
+ bl_int_37_13 bl_int_36_13 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c14
+ bl_int_37_14 bl_int_36_14 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c15
+ bl_int_37_15 bl_int_36_15 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c16
+ bl_int_37_16 bl_int_36_16 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c17
+ bl_int_37_17 bl_int_36_17 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c18
+ bl_int_37_18 bl_int_36_18 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c19
+ bl_int_37_19 bl_int_36_19 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c20
+ bl_int_37_20 bl_int_36_20 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c21
+ bl_int_37_21 bl_int_36_21 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c22
+ bl_int_37_22 bl_int_36_22 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c23
+ bl_int_37_23 bl_int_36_23 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c24
+ bl_int_37_24 bl_int_36_24 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c25
+ bl_int_37_25 bl_int_36_25 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c26
+ bl_int_37_26 bl_int_36_26 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c27
+ bl_int_37_27 bl_int_36_27 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c28
+ bl_int_37_28 bl_int_36_28 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c29
+ bl_int_37_29 bl_int_36_29 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c30
+ bl_int_37_30 bl_int_36_30 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c31
+ bl_int_37_31 bl_int_36_31 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c32
+ bl_int_37_32 bl_int_36_32 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c33
+ bl_int_37_33 bl_int_36_33 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c34
+ bl_int_37_34 bl_int_36_34 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c35
+ bl_int_37_35 bl_int_36_35 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c36
+ bl_int_37_36 bl_int_36_36 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c37
+ bl_int_37_37 bl_int_36_37 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c38
+ bl_int_37_38 bl_int_36_38 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c39
+ bl_int_37_39 bl_int_36_39 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c40
+ bl_int_37_40 bl_int_36_40 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c41
+ bl_int_37_41 bl_int_36_41 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c42
+ bl_int_37_42 bl_int_36_42 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c43
+ bl_int_37_43 bl_int_36_43 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c44
+ bl_int_37_44 bl_int_36_44 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c45
+ bl_int_37_45 bl_int_36_45 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c46
+ bl_int_37_46 bl_int_36_46 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c47
+ bl_int_37_47 bl_int_36_47 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c48
+ bl_int_37_48 bl_int_36_48 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c49
+ bl_int_37_49 bl_int_36_49 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c50
+ bl_int_37_50 bl_int_36_50 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c51
+ bl_int_37_51 bl_int_36_51 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c52
+ bl_int_37_52 bl_int_36_52 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c53
+ bl_int_37_53 bl_int_36_53 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c54
+ bl_int_37_54 bl_int_36_54 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c55
+ bl_int_37_55 bl_int_36_55 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c56
+ bl_int_37_56 bl_int_36_56 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c57
+ bl_int_37_57 bl_int_36_57 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c58
+ bl_int_37_58 bl_int_36_58 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c59
+ bl_int_37_59 bl_int_36_59 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c60
+ bl_int_37_60 bl_int_36_60 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c61
+ bl_int_37_61 bl_int_36_61 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c62
+ bl_int_37_62 bl_int_36_62 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c63
+ bl_int_37_63 bl_int_36_63 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c64
+ bl_int_37_64 bl_int_36_64 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c65
+ bl_int_37_65 bl_int_36_65 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c66
+ bl_int_37_66 bl_int_36_66 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c67
+ bl_int_37_67 bl_int_36_67 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c68
+ bl_int_37_68 bl_int_36_68 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c69
+ bl_int_37_69 bl_int_36_69 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c70
+ bl_int_37_70 bl_int_36_70 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c71
+ bl_int_37_71 bl_int_36_71 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c72
+ bl_int_37_72 bl_int_36_72 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c73
+ bl_int_37_73 bl_int_36_73 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c74
+ bl_int_37_74 bl_int_36_74 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c75
+ bl_int_37_75 bl_int_36_75 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c76
+ bl_int_37_76 bl_int_36_76 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c77
+ bl_int_37_77 bl_int_36_77 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c78
+ bl_int_37_78 bl_int_36_78 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c79
+ bl_int_37_79 bl_int_36_79 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c80
+ bl_int_37_80 bl_int_36_80 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c81
+ bl_int_37_81 bl_int_36_81 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c82
+ bl_int_37_82 bl_int_36_82 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c83
+ bl_int_37_83 bl_int_36_83 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c84
+ bl_int_37_84 bl_int_36_84 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c85
+ bl_int_37_85 bl_int_36_85 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c86
+ bl_int_37_86 bl_int_36_86 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c87
+ bl_int_37_87 bl_int_36_87 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c88
+ bl_int_37_88 bl_int_36_88 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c89
+ bl_int_37_89 bl_int_36_89 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c90
+ bl_int_37_90 bl_int_36_90 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c91
+ bl_int_37_91 bl_int_36_91 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c92
+ bl_int_37_92 bl_int_36_92 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c93
+ bl_int_37_93 bl_int_36_93 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c94
+ bl_int_37_94 bl_int_36_94 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c95
+ bl_int_37_95 bl_int_36_95 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c96
+ bl_int_37_96 bl_int_36_96 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c97
+ bl_int_37_97 bl_int_36_97 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c98
+ bl_int_37_98 bl_int_36_98 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c99
+ bl_int_37_99 bl_int_36_99 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c100
+ bl_int_37_100 bl_int_36_100 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c101
+ bl_int_37_101 bl_int_36_101 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c102
+ bl_int_37_102 bl_int_36_102 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c103
+ bl_int_37_103 bl_int_36_103 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c104
+ bl_int_37_104 bl_int_36_104 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c105
+ bl_int_37_105 bl_int_36_105 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c106
+ bl_int_37_106 bl_int_36_106 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c107
+ bl_int_37_107 bl_int_36_107 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c108
+ bl_int_37_108 bl_int_36_108 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c109
+ bl_int_37_109 bl_int_36_109 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c110
+ bl_int_37_110 bl_int_36_110 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c111
+ bl_int_37_111 bl_int_36_111 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c112
+ bl_int_37_112 bl_int_36_112 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c113
+ bl_int_37_113 bl_int_36_113 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c114
+ bl_int_37_114 bl_int_36_114 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c115
+ bl_int_37_115 bl_int_36_115 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c116
+ bl_int_37_116 bl_int_36_116 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c117
+ bl_int_37_117 bl_int_36_117 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c118
+ bl_int_37_118 bl_int_36_118 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c119
+ bl_int_37_119 bl_int_36_119 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c120
+ bl_int_37_120 bl_int_36_120 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c121
+ bl_int_37_121 bl_int_36_121 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c122
+ bl_int_37_122 bl_int_36_122 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c123
+ bl_int_37_123 bl_int_36_123 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c124
+ bl_int_37_124 bl_int_36_124 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c125
+ bl_int_37_125 bl_int_36_125 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c126
+ bl_int_37_126 bl_int_36_126 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c127
+ bl_int_37_127 bl_int_36_127 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c128
+ bl_int_37_128 bl_int_36_128 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c129
+ bl_int_37_129 bl_int_36_129 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c130
+ bl_int_37_130 bl_int_36_130 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c131
+ bl_int_37_131 bl_int_36_131 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c132
+ bl_int_37_132 bl_int_36_132 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c133
+ bl_int_37_133 bl_int_36_133 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c134
+ bl_int_37_134 bl_int_36_134 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c135
+ bl_int_37_135 bl_int_36_135 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c136
+ bl_int_37_136 bl_int_36_136 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c137
+ bl_int_37_137 bl_int_36_137 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c138
+ bl_int_37_138 bl_int_36_138 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c139
+ bl_int_37_139 bl_int_36_139 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c140
+ bl_int_37_140 bl_int_36_140 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c141
+ bl_int_37_141 bl_int_36_141 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c142
+ bl_int_37_142 bl_int_36_142 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c143
+ bl_int_37_143 bl_int_36_143 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c144
+ bl_int_37_144 bl_int_36_144 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c145
+ bl_int_37_145 bl_int_36_145 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c146
+ bl_int_37_146 bl_int_36_146 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c147
+ bl_int_37_147 bl_int_36_147 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c148
+ bl_int_37_148 bl_int_36_148 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c149
+ bl_int_37_149 bl_int_36_149 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c150
+ bl_int_37_150 bl_int_36_150 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c151
+ bl_int_37_151 bl_int_36_151 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c152
+ bl_int_37_152 bl_int_36_152 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c153
+ bl_int_37_153 bl_int_36_153 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c154
+ bl_int_37_154 bl_int_36_154 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c155
+ bl_int_37_155 bl_int_36_155 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c156
+ bl_int_37_156 bl_int_36_156 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c157
+ bl_int_37_157 bl_int_36_157 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c158
+ bl_int_37_158 bl_int_36_158 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c159
+ bl_int_37_159 bl_int_36_159 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c160
+ bl_int_37_160 bl_int_36_160 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c161
+ bl_int_37_161 bl_int_36_161 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c162
+ bl_int_37_162 bl_int_36_162 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c163
+ bl_int_37_163 bl_int_36_163 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c164
+ bl_int_37_164 bl_int_36_164 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c165
+ bl_int_37_165 bl_int_36_165 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c166
+ bl_int_37_166 bl_int_36_166 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c167
+ bl_int_37_167 bl_int_36_167 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c168
+ bl_int_37_168 bl_int_36_168 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c169
+ bl_int_37_169 bl_int_36_169 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c170
+ bl_int_37_170 bl_int_36_170 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c171
+ bl_int_37_171 bl_int_36_171 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c172
+ bl_int_37_172 bl_int_36_172 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c173
+ bl_int_37_173 bl_int_36_173 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c174
+ bl_int_37_174 bl_int_36_174 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c175
+ bl_int_37_175 bl_int_36_175 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c176
+ bl_int_37_176 bl_int_36_176 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c177
+ bl_int_37_177 bl_int_36_177 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c178
+ bl_int_37_178 bl_int_36_178 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c179
+ bl_int_37_179 bl_int_36_179 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c180
+ bl_int_37_180 bl_int_36_180 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c181
+ bl_int_37_181 bl_int_36_181 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c182
+ bl_int_37_182 bl_int_36_182 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r37_c183
+ bl_int_37_183 bl_int_36_183 wl_0_37 gnd
+ sram_rom_base_one_cell
Xbit_r38_c0
+ bl_int_38_0 bl_int_37_0 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c1
+ bl_int_38_1 bl_int_37_1 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c2
+ bl_int_38_2 bl_int_37_2 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c3
+ bl_int_38_3 bl_int_37_3 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c4
+ bl_int_38_4 bl_int_37_4 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c5
+ bl_int_38_5 bl_int_37_5 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c6
+ bl_int_38_6 bl_int_37_6 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c7
+ bl_int_38_7 bl_int_37_7 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c8
+ bl_int_38_8 bl_int_37_8 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c9
+ bl_int_38_9 bl_int_37_9 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c10
+ bl_int_38_10 bl_int_37_10 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c11
+ bl_int_38_11 bl_int_37_11 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c12
+ bl_int_38_12 bl_int_37_12 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c13
+ bl_int_38_13 bl_int_37_13 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c14
+ bl_int_38_14 bl_int_37_14 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c15
+ bl_int_38_15 bl_int_37_15 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c16
+ bl_int_38_16 bl_int_37_16 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c17
+ bl_int_38_17 bl_int_37_17 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c18
+ bl_int_38_18 bl_int_37_18 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c19
+ bl_int_38_19 bl_int_37_19 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c20
+ bl_int_38_20 bl_int_37_20 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c21
+ bl_int_38_21 bl_int_37_21 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c22
+ bl_int_38_22 bl_int_37_22 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c23
+ bl_int_38_23 bl_int_37_23 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c24
+ bl_int_38_24 bl_int_37_24 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c25
+ bl_int_38_25 bl_int_37_25 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c26
+ bl_int_38_26 bl_int_37_26 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c27
+ bl_int_38_27 bl_int_37_27 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c28
+ bl_int_38_28 bl_int_37_28 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c29
+ bl_int_38_29 bl_int_37_29 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c30
+ bl_int_38_30 bl_int_37_30 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c31
+ bl_int_38_31 bl_int_37_31 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c32
+ bl_int_38_32 bl_int_37_32 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c33
+ bl_int_38_33 bl_int_37_33 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c34
+ bl_int_38_34 bl_int_37_34 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c35
+ bl_int_38_35 bl_int_37_35 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c36
+ bl_int_38_36 bl_int_37_36 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c37
+ bl_int_38_37 bl_int_37_37 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c38
+ bl_int_38_38 bl_int_37_38 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c39
+ bl_int_38_39 bl_int_37_39 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c40
+ bl_int_38_40 bl_int_37_40 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c41
+ bl_int_38_41 bl_int_37_41 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c42
+ bl_int_38_42 bl_int_37_42 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c43
+ bl_int_38_43 bl_int_37_43 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c44
+ bl_int_38_44 bl_int_37_44 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c45
+ bl_int_38_45 bl_int_37_45 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c46
+ bl_int_38_46 bl_int_37_46 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c47
+ bl_int_38_47 bl_int_37_47 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c48
+ bl_int_38_48 bl_int_37_48 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c49
+ bl_int_38_49 bl_int_37_49 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c50
+ bl_int_38_50 bl_int_37_50 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c51
+ bl_int_38_51 bl_int_37_51 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c52
+ bl_int_38_52 bl_int_37_52 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c53
+ bl_int_38_53 bl_int_37_53 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c54
+ bl_int_38_54 bl_int_37_54 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c55
+ bl_int_38_55 bl_int_37_55 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c56
+ bl_int_38_56 bl_int_37_56 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c57
+ bl_int_38_57 bl_int_37_57 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c58
+ bl_int_38_58 bl_int_37_58 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c59
+ bl_int_38_59 bl_int_37_59 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c60
+ bl_int_38_60 bl_int_37_60 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c61
+ bl_int_38_61 bl_int_37_61 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c62
+ bl_int_38_62 bl_int_37_62 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c63
+ bl_int_38_63 bl_int_37_63 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c64
+ bl_int_38_64 bl_int_37_64 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c65
+ bl_int_38_65 bl_int_37_65 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c66
+ bl_int_38_66 bl_int_37_66 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c67
+ bl_int_38_67 bl_int_37_67 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c68
+ bl_int_38_68 bl_int_37_68 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c69
+ bl_int_38_69 bl_int_37_69 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c70
+ bl_int_38_70 bl_int_37_70 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c71
+ bl_int_38_71 bl_int_37_71 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c72
+ bl_int_38_72 bl_int_37_72 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c73
+ bl_int_38_73 bl_int_37_73 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c74
+ bl_int_38_74 bl_int_37_74 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c75
+ bl_int_38_75 bl_int_37_75 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c76
+ bl_int_38_76 bl_int_37_76 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c77
+ bl_int_38_77 bl_int_37_77 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c78
+ bl_int_38_78 bl_int_37_78 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c79
+ bl_int_38_79 bl_int_37_79 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c80
+ bl_int_38_80 bl_int_37_80 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c81
+ bl_int_38_81 bl_int_37_81 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c82
+ bl_int_38_82 bl_int_37_82 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c83
+ bl_int_38_83 bl_int_37_83 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c84
+ bl_int_38_84 bl_int_37_84 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c85
+ bl_int_38_85 bl_int_37_85 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c86
+ bl_int_38_86 bl_int_37_86 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c87
+ bl_int_38_87 bl_int_37_87 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c88
+ bl_int_38_88 bl_int_37_88 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c89
+ bl_int_38_89 bl_int_37_89 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c90
+ bl_int_38_90 bl_int_37_90 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c91
+ bl_int_38_91 bl_int_37_91 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c92
+ bl_int_38_92 bl_int_37_92 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c93
+ bl_int_38_93 bl_int_37_93 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c94
+ bl_int_38_94 bl_int_37_94 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c95
+ bl_int_38_95 bl_int_37_95 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c96
+ bl_int_38_96 bl_int_37_96 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c97
+ bl_int_38_97 bl_int_37_97 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c98
+ bl_int_38_98 bl_int_37_98 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c99
+ bl_int_38_99 bl_int_37_99 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c100
+ bl_int_38_100 bl_int_37_100 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c101
+ bl_int_38_101 bl_int_37_101 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c102
+ bl_int_38_102 bl_int_37_102 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c103
+ bl_int_38_103 bl_int_37_103 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c104
+ bl_int_38_104 bl_int_37_104 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c105
+ bl_int_38_105 bl_int_37_105 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c106
+ bl_int_38_106 bl_int_37_106 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c107
+ bl_int_38_107 bl_int_37_107 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c108
+ bl_int_38_108 bl_int_37_108 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c109
+ bl_int_38_109 bl_int_37_109 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c110
+ bl_int_38_110 bl_int_37_110 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c111
+ bl_int_38_111 bl_int_37_111 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c112
+ bl_int_38_112 bl_int_37_112 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c113
+ bl_int_38_113 bl_int_37_113 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c114
+ bl_int_38_114 bl_int_37_114 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c115
+ bl_int_38_115 bl_int_37_115 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c116
+ bl_int_38_116 bl_int_37_116 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c117
+ bl_int_38_117 bl_int_37_117 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c118
+ bl_int_38_118 bl_int_37_118 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c119
+ bl_int_38_119 bl_int_37_119 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c120
+ bl_int_38_120 bl_int_37_120 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c121
+ bl_int_38_121 bl_int_37_121 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c122
+ bl_int_38_122 bl_int_37_122 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c123
+ bl_int_38_123 bl_int_37_123 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c124
+ bl_int_38_124 bl_int_37_124 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c125
+ bl_int_38_125 bl_int_37_125 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c126
+ bl_int_38_126 bl_int_37_126 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c127
+ bl_int_38_127 bl_int_37_127 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c128
+ bl_int_38_128 bl_int_37_128 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c129
+ bl_int_38_129 bl_int_37_129 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c130
+ bl_int_38_130 bl_int_37_130 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c131
+ bl_int_38_131 bl_int_37_131 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c132
+ bl_int_38_132 bl_int_37_132 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c133
+ bl_int_38_133 bl_int_37_133 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c134
+ bl_int_38_134 bl_int_37_134 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c135
+ bl_int_38_135 bl_int_37_135 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c136
+ bl_int_38_136 bl_int_37_136 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c137
+ bl_int_38_137 bl_int_37_137 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c138
+ bl_int_38_138 bl_int_37_138 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c139
+ bl_int_38_139 bl_int_37_139 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c140
+ bl_int_38_140 bl_int_37_140 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c141
+ bl_int_38_141 bl_int_37_141 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c142
+ bl_int_38_142 bl_int_37_142 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c143
+ bl_int_38_143 bl_int_37_143 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c144
+ bl_int_38_144 bl_int_37_144 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c145
+ bl_int_38_145 bl_int_37_145 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c146
+ bl_int_38_146 bl_int_37_146 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c147
+ bl_int_38_147 bl_int_37_147 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c148
+ bl_int_38_148 bl_int_37_148 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c149
+ bl_int_38_149 bl_int_37_149 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c150
+ bl_int_38_150 bl_int_37_150 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c151
+ bl_int_38_151 bl_int_37_151 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c152
+ bl_int_38_152 bl_int_37_152 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c153
+ bl_int_38_153 bl_int_37_153 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c154
+ bl_int_38_154 bl_int_37_154 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c155
+ bl_int_38_155 bl_int_37_155 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c156
+ bl_int_38_156 bl_int_37_156 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c157
+ bl_int_38_157 bl_int_37_157 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c158
+ bl_int_38_158 bl_int_37_158 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c159
+ bl_int_38_159 bl_int_37_159 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c160
+ bl_int_38_160 bl_int_37_160 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c161
+ bl_int_38_161 bl_int_37_161 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c162
+ bl_int_38_162 bl_int_37_162 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c163
+ bl_int_38_163 bl_int_37_163 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c164
+ bl_int_38_164 bl_int_37_164 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c165
+ bl_int_38_165 bl_int_37_165 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c166
+ bl_int_38_166 bl_int_37_166 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c167
+ bl_int_38_167 bl_int_37_167 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c168
+ bl_int_38_168 bl_int_37_168 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c169
+ bl_int_38_169 bl_int_37_169 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c170
+ bl_int_38_170 bl_int_37_170 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c171
+ bl_int_38_171 bl_int_37_171 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c172
+ bl_int_38_172 bl_int_37_172 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c173
+ bl_int_38_173 bl_int_37_173 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c174
+ bl_int_38_174 bl_int_37_174 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c175
+ bl_int_38_175 bl_int_37_175 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c176
+ bl_int_38_176 bl_int_37_176 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c177
+ bl_int_38_177 bl_int_37_177 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c178
+ bl_int_38_178 bl_int_37_178 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c179
+ bl_int_38_179 bl_int_37_179 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c180
+ bl_int_38_180 bl_int_37_180 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c181
+ bl_int_38_181 bl_int_37_181 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c182
+ bl_int_38_182 bl_int_37_182 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r38_c183
+ bl_int_38_183 bl_int_37_183 wl_0_38 gnd
+ sram_rom_base_one_cell
Xbit_r39_c0
+ bl_int_39_0 bl_int_38_0 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c1
+ bl_int_39_1 bl_int_38_1 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c2
+ bl_int_39_2 bl_int_38_2 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c3
+ bl_int_39_3 bl_int_38_3 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c4
+ bl_int_39_4 bl_int_38_4 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c5
+ bl_int_39_5 bl_int_38_5 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c6
+ bl_int_39_6 bl_int_38_6 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c7
+ bl_int_39_7 bl_int_38_7 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c8
+ bl_int_39_8 bl_int_38_8 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c9
+ bl_int_39_9 bl_int_38_9 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c10
+ bl_int_39_10 bl_int_38_10 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c11
+ bl_int_39_11 bl_int_38_11 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c12
+ bl_int_39_12 bl_int_38_12 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c13
+ bl_int_39_13 bl_int_38_13 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c14
+ bl_int_39_14 bl_int_38_14 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c15
+ bl_int_39_15 bl_int_38_15 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c16
+ bl_int_39_16 bl_int_38_16 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c17
+ bl_int_39_17 bl_int_38_17 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c18
+ bl_int_39_18 bl_int_38_18 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c19
+ bl_int_39_19 bl_int_38_19 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c20
+ bl_int_39_20 bl_int_38_20 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c21
+ bl_int_39_21 bl_int_38_21 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c22
+ bl_int_39_22 bl_int_38_22 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c23
+ bl_int_39_23 bl_int_38_23 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c24
+ bl_int_39_24 bl_int_38_24 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c25
+ bl_int_39_25 bl_int_38_25 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c26
+ bl_int_39_26 bl_int_38_26 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c27
+ bl_int_39_27 bl_int_38_27 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c28
+ bl_int_39_28 bl_int_38_28 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c29
+ bl_int_39_29 bl_int_38_29 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c30
+ bl_int_39_30 bl_int_38_30 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c31
+ bl_int_39_31 bl_int_38_31 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c32
+ bl_int_39_32 bl_int_38_32 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c33
+ bl_int_39_33 bl_int_38_33 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c34
+ bl_int_39_34 bl_int_38_34 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c35
+ bl_int_39_35 bl_int_38_35 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c36
+ bl_int_39_36 bl_int_38_36 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c37
+ bl_int_39_37 bl_int_38_37 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c38
+ bl_int_39_38 bl_int_38_38 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c39
+ bl_int_39_39 bl_int_38_39 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c40
+ bl_int_39_40 bl_int_38_40 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c41
+ bl_int_39_41 bl_int_38_41 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c42
+ bl_int_39_42 bl_int_38_42 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c43
+ bl_int_39_43 bl_int_38_43 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c44
+ bl_int_39_44 bl_int_38_44 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c45
+ bl_int_39_45 bl_int_38_45 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c46
+ bl_int_39_46 bl_int_38_46 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c47
+ bl_int_39_47 bl_int_38_47 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c48
+ bl_int_39_48 bl_int_38_48 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c49
+ bl_int_39_49 bl_int_38_49 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c50
+ bl_int_39_50 bl_int_38_50 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c51
+ bl_int_39_51 bl_int_38_51 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c52
+ bl_int_39_52 bl_int_38_52 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c53
+ bl_int_39_53 bl_int_38_53 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c54
+ bl_int_39_54 bl_int_38_54 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c55
+ bl_int_39_55 bl_int_38_55 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c56
+ bl_int_39_56 bl_int_38_56 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c57
+ bl_int_39_57 bl_int_38_57 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c58
+ bl_int_39_58 bl_int_38_58 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c59
+ bl_int_39_59 bl_int_38_59 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c60
+ bl_int_39_60 bl_int_38_60 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c61
+ bl_int_39_61 bl_int_38_61 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c62
+ bl_int_39_62 bl_int_38_62 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c63
+ bl_int_39_63 bl_int_38_63 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c64
+ bl_int_39_64 bl_int_38_64 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c65
+ bl_int_39_65 bl_int_38_65 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c66
+ bl_int_39_66 bl_int_38_66 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c67
+ bl_int_39_67 bl_int_38_67 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c68
+ bl_int_39_68 bl_int_38_68 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c69
+ bl_int_39_69 bl_int_38_69 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c70
+ bl_int_39_70 bl_int_38_70 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c71
+ bl_int_39_71 bl_int_38_71 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c72
+ bl_int_39_72 bl_int_38_72 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c73
+ bl_int_39_73 bl_int_38_73 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c74
+ bl_int_39_74 bl_int_38_74 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c75
+ bl_int_39_75 bl_int_38_75 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c76
+ bl_int_39_76 bl_int_38_76 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c77
+ bl_int_39_77 bl_int_38_77 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c78
+ bl_int_39_78 bl_int_38_78 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c79
+ bl_int_39_79 bl_int_38_79 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c80
+ bl_int_39_80 bl_int_38_80 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c81
+ bl_int_39_81 bl_int_38_81 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c82
+ bl_int_39_82 bl_int_38_82 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c83
+ bl_int_39_83 bl_int_38_83 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c84
+ bl_int_39_84 bl_int_38_84 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c85
+ bl_int_39_85 bl_int_38_85 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c86
+ bl_int_39_86 bl_int_38_86 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c87
+ bl_int_39_87 bl_int_38_87 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c88
+ bl_int_39_88 bl_int_38_88 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c89
+ bl_int_39_89 bl_int_38_89 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c90
+ bl_int_39_90 bl_int_38_90 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c91
+ bl_int_39_91 bl_int_38_91 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c92
+ bl_int_39_92 bl_int_38_92 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c93
+ bl_int_39_93 bl_int_38_93 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c94
+ bl_int_39_94 bl_int_38_94 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c95
+ bl_int_39_95 bl_int_38_95 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c96
+ bl_int_39_96 bl_int_38_96 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c97
+ bl_int_39_97 bl_int_38_97 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c98
+ bl_int_39_98 bl_int_38_98 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c99
+ bl_int_39_99 bl_int_38_99 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c100
+ bl_int_39_100 bl_int_38_100 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c101
+ bl_int_39_101 bl_int_38_101 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c102
+ bl_int_39_102 bl_int_38_102 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c103
+ bl_int_39_103 bl_int_38_103 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c104
+ bl_int_39_104 bl_int_38_104 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c105
+ bl_int_39_105 bl_int_38_105 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c106
+ bl_int_39_106 bl_int_38_106 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c107
+ bl_int_39_107 bl_int_38_107 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c108
+ bl_int_39_108 bl_int_38_108 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c109
+ bl_int_39_109 bl_int_38_109 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c110
+ bl_int_39_110 bl_int_38_110 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c111
+ bl_int_39_111 bl_int_38_111 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c112
+ bl_int_39_112 bl_int_38_112 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c113
+ bl_int_39_113 bl_int_38_113 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c114
+ bl_int_39_114 bl_int_38_114 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c115
+ bl_int_39_115 bl_int_38_115 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c116
+ bl_int_39_116 bl_int_38_116 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c117
+ bl_int_39_117 bl_int_38_117 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c118
+ bl_int_39_118 bl_int_38_118 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c119
+ bl_int_39_119 bl_int_38_119 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c120
+ bl_int_39_120 bl_int_38_120 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c121
+ bl_int_39_121 bl_int_38_121 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c122
+ bl_int_39_122 bl_int_38_122 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c123
+ bl_int_39_123 bl_int_38_123 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c124
+ bl_int_39_124 bl_int_38_124 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c125
+ bl_int_39_125 bl_int_38_125 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c126
+ bl_int_39_126 bl_int_38_126 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c127
+ bl_int_39_127 bl_int_38_127 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c128
+ bl_int_39_128 bl_int_38_128 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c129
+ bl_int_39_129 bl_int_38_129 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c130
+ bl_int_39_130 bl_int_38_130 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c131
+ bl_int_39_131 bl_int_38_131 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c132
+ bl_int_39_132 bl_int_38_132 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c133
+ bl_int_39_133 bl_int_38_133 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c134
+ bl_int_39_134 bl_int_38_134 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c135
+ bl_int_39_135 bl_int_38_135 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c136
+ bl_int_39_136 bl_int_38_136 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c137
+ bl_int_39_137 bl_int_38_137 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c138
+ bl_int_39_138 bl_int_38_138 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c139
+ bl_int_39_139 bl_int_38_139 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c140
+ bl_int_39_140 bl_int_38_140 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c141
+ bl_int_39_141 bl_int_38_141 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c142
+ bl_int_39_142 bl_int_38_142 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c143
+ bl_int_39_143 bl_int_38_143 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c144
+ bl_int_39_144 bl_int_38_144 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c145
+ bl_int_39_145 bl_int_38_145 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c146
+ bl_int_39_146 bl_int_38_146 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c147
+ bl_int_39_147 bl_int_38_147 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c148
+ bl_int_39_148 bl_int_38_148 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c149
+ bl_int_39_149 bl_int_38_149 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c150
+ bl_int_39_150 bl_int_38_150 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c151
+ bl_int_39_151 bl_int_38_151 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c152
+ bl_int_39_152 bl_int_38_152 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c153
+ bl_int_39_153 bl_int_38_153 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c154
+ bl_int_39_154 bl_int_38_154 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c155
+ bl_int_39_155 bl_int_38_155 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c156
+ bl_int_39_156 bl_int_38_156 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c157
+ bl_int_39_157 bl_int_38_157 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c158
+ bl_int_39_158 bl_int_38_158 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c159
+ bl_int_39_159 bl_int_38_159 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c160
+ bl_int_39_160 bl_int_38_160 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c161
+ bl_int_39_161 bl_int_38_161 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c162
+ bl_int_39_162 bl_int_38_162 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c163
+ bl_int_39_163 bl_int_38_163 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c164
+ bl_int_39_164 bl_int_38_164 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c165
+ bl_int_39_165 bl_int_38_165 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c166
+ bl_int_39_166 bl_int_38_166 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c167
+ bl_int_39_167 bl_int_38_167 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c168
+ bl_int_39_168 bl_int_38_168 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c169
+ bl_int_39_169 bl_int_38_169 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c170
+ bl_int_39_170 bl_int_38_170 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c171
+ bl_int_39_171 bl_int_38_171 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c172
+ bl_int_39_172 bl_int_38_172 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c173
+ bl_int_39_173 bl_int_38_173 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c174
+ bl_int_39_174 bl_int_38_174 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c175
+ bl_int_39_175 bl_int_38_175 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c176
+ bl_int_39_176 bl_int_38_176 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c177
+ bl_int_39_177 bl_int_38_177 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c178
+ bl_int_39_178 bl_int_38_178 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c179
+ bl_int_39_179 bl_int_38_179 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c180
+ bl_int_39_180 bl_int_38_180 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c181
+ bl_int_39_181 bl_int_38_181 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c182
+ bl_int_39_182 bl_int_38_182 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r39_c183
+ bl_int_39_183 bl_int_38_183 wl_0_39 gnd
+ sram_rom_base_one_cell
Xbit_r40_c0
+ bl_int_40_0 bl_int_39_0 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c1
+ bl_int_40_1 bl_int_39_1 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c2
+ bl_int_40_2 bl_int_39_2 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c3
+ bl_int_40_3 bl_int_39_3 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c4
+ bl_int_40_4 bl_int_39_4 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c5
+ bl_int_40_5 bl_int_39_5 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c6
+ bl_int_40_6 bl_int_39_6 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c7
+ bl_int_40_7 bl_int_39_7 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c8
+ bl_int_40_8 bl_int_39_8 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c9
+ bl_int_40_9 bl_int_39_9 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c10
+ bl_int_40_10 bl_int_39_10 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c11
+ bl_int_40_11 bl_int_39_11 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c12
+ bl_int_40_12 bl_int_39_12 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c13
+ bl_int_40_13 bl_int_39_13 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c14
+ bl_int_40_14 bl_int_39_14 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c15
+ bl_int_40_15 bl_int_39_15 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c16
+ bl_int_40_16 bl_int_39_16 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c17
+ bl_int_40_17 bl_int_39_17 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c18
+ bl_int_40_18 bl_int_39_18 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c19
+ bl_int_40_19 bl_int_39_19 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c20
+ bl_int_40_20 bl_int_39_20 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c21
+ bl_int_40_21 bl_int_39_21 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c22
+ bl_int_40_22 bl_int_39_22 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c23
+ bl_int_40_23 bl_int_39_23 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c24
+ bl_int_40_24 bl_int_39_24 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c25
+ bl_int_40_25 bl_int_39_25 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c26
+ bl_int_40_26 bl_int_39_26 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c27
+ bl_int_40_27 bl_int_39_27 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c28
+ bl_int_40_28 bl_int_39_28 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c29
+ bl_int_40_29 bl_int_39_29 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c30
+ bl_int_40_30 bl_int_39_30 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c31
+ bl_int_40_31 bl_int_39_31 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c32
+ bl_int_40_32 bl_int_39_32 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c33
+ bl_int_40_33 bl_int_39_33 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c34
+ bl_int_40_34 bl_int_39_34 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c35
+ bl_int_40_35 bl_int_39_35 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c36
+ bl_int_40_36 bl_int_39_36 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c37
+ bl_int_40_37 bl_int_39_37 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c38
+ bl_int_40_38 bl_int_39_38 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c39
+ bl_int_40_39 bl_int_39_39 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c40
+ bl_int_40_40 bl_int_39_40 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c41
+ bl_int_40_41 bl_int_39_41 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c42
+ bl_int_40_42 bl_int_39_42 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c43
+ bl_int_40_43 bl_int_39_43 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c44
+ bl_int_40_44 bl_int_39_44 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c45
+ bl_int_40_45 bl_int_39_45 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c46
+ bl_int_40_46 bl_int_39_46 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c47
+ bl_int_40_47 bl_int_39_47 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c48
+ bl_int_40_48 bl_int_39_48 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c49
+ bl_int_40_49 bl_int_39_49 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c50
+ bl_int_40_50 bl_int_39_50 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c51
+ bl_int_40_51 bl_int_39_51 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c52
+ bl_int_40_52 bl_int_39_52 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c53
+ bl_int_40_53 bl_int_39_53 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c54
+ bl_int_40_54 bl_int_39_54 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c55
+ bl_int_40_55 bl_int_39_55 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c56
+ bl_int_40_56 bl_int_39_56 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c57
+ bl_int_40_57 bl_int_39_57 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c58
+ bl_int_40_58 bl_int_39_58 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c59
+ bl_int_40_59 bl_int_39_59 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c60
+ bl_int_40_60 bl_int_39_60 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c61
+ bl_int_40_61 bl_int_39_61 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c62
+ bl_int_40_62 bl_int_39_62 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c63
+ bl_int_40_63 bl_int_39_63 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c64
+ bl_int_40_64 bl_int_39_64 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c65
+ bl_int_40_65 bl_int_39_65 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c66
+ bl_int_40_66 bl_int_39_66 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c67
+ bl_int_40_67 bl_int_39_67 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c68
+ bl_int_40_68 bl_int_39_68 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c69
+ bl_int_40_69 bl_int_39_69 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c70
+ bl_int_40_70 bl_int_39_70 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c71
+ bl_int_40_71 bl_int_39_71 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c72
+ bl_int_40_72 bl_int_39_72 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c73
+ bl_int_40_73 bl_int_39_73 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c74
+ bl_int_40_74 bl_int_39_74 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c75
+ bl_int_40_75 bl_int_39_75 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c76
+ bl_int_40_76 bl_int_39_76 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c77
+ bl_int_40_77 bl_int_39_77 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c78
+ bl_int_40_78 bl_int_39_78 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c79
+ bl_int_40_79 bl_int_39_79 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c80
+ bl_int_40_80 bl_int_39_80 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c81
+ bl_int_40_81 bl_int_39_81 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c82
+ bl_int_40_82 bl_int_39_82 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c83
+ bl_int_40_83 bl_int_39_83 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c84
+ bl_int_40_84 bl_int_39_84 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c85
+ bl_int_40_85 bl_int_39_85 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c86
+ bl_int_40_86 bl_int_39_86 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c87
+ bl_int_40_87 bl_int_39_87 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c88
+ bl_int_40_88 bl_int_39_88 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c89
+ bl_int_40_89 bl_int_39_89 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c90
+ bl_int_40_90 bl_int_39_90 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c91
+ bl_int_40_91 bl_int_39_91 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c92
+ bl_int_40_92 bl_int_39_92 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c93
+ bl_int_40_93 bl_int_39_93 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c94
+ bl_int_40_94 bl_int_39_94 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c95
+ bl_int_40_95 bl_int_39_95 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c96
+ bl_int_40_96 bl_int_39_96 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c97
+ bl_int_40_97 bl_int_39_97 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c98
+ bl_int_40_98 bl_int_39_98 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c99
+ bl_int_40_99 bl_int_39_99 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c100
+ bl_int_40_100 bl_int_39_100 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c101
+ bl_int_40_101 bl_int_39_101 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c102
+ bl_int_40_102 bl_int_39_102 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c103
+ bl_int_40_103 bl_int_39_103 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c104
+ bl_int_40_104 bl_int_39_104 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c105
+ bl_int_40_105 bl_int_39_105 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c106
+ bl_int_40_106 bl_int_39_106 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c107
+ bl_int_40_107 bl_int_39_107 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c108
+ bl_int_40_108 bl_int_39_108 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c109
+ bl_int_40_109 bl_int_39_109 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c110
+ bl_int_40_110 bl_int_39_110 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c111
+ bl_int_40_111 bl_int_39_111 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c112
+ bl_int_40_112 bl_int_39_112 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c113
+ bl_int_40_113 bl_int_39_113 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c114
+ bl_int_40_114 bl_int_39_114 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c115
+ bl_int_40_115 bl_int_39_115 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c116
+ bl_int_40_116 bl_int_39_116 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c117
+ bl_int_40_117 bl_int_39_117 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c118
+ bl_int_40_118 bl_int_39_118 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c119
+ bl_int_40_119 bl_int_39_119 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c120
+ bl_int_40_120 bl_int_39_120 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c121
+ bl_int_40_121 bl_int_39_121 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c122
+ bl_int_40_122 bl_int_39_122 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c123
+ bl_int_40_123 bl_int_39_123 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c124
+ bl_int_40_124 bl_int_39_124 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c125
+ bl_int_40_125 bl_int_39_125 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c126
+ bl_int_40_126 bl_int_39_126 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c127
+ bl_int_40_127 bl_int_39_127 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c128
+ bl_int_40_128 bl_int_39_128 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c129
+ bl_int_40_129 bl_int_39_129 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c130
+ bl_int_40_130 bl_int_39_130 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c131
+ bl_int_40_131 bl_int_39_131 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c132
+ bl_int_40_132 bl_int_39_132 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c133
+ bl_int_40_133 bl_int_39_133 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c134
+ bl_int_40_134 bl_int_39_134 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c135
+ bl_int_40_135 bl_int_39_135 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c136
+ bl_int_40_136 bl_int_39_136 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c137
+ bl_int_40_137 bl_int_39_137 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c138
+ bl_int_40_138 bl_int_39_138 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c139
+ bl_int_40_139 bl_int_39_139 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c140
+ bl_int_40_140 bl_int_39_140 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c141
+ bl_int_40_141 bl_int_39_141 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c142
+ bl_int_40_142 bl_int_39_142 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c143
+ bl_int_40_143 bl_int_39_143 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c144
+ bl_int_40_144 bl_int_39_144 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c145
+ bl_int_40_145 bl_int_39_145 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c146
+ bl_int_40_146 bl_int_39_146 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c147
+ bl_int_40_147 bl_int_39_147 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c148
+ bl_int_40_148 bl_int_39_148 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c149
+ bl_int_40_149 bl_int_39_149 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c150
+ bl_int_40_150 bl_int_39_150 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c151
+ bl_int_40_151 bl_int_39_151 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c152
+ bl_int_40_152 bl_int_39_152 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c153
+ bl_int_40_153 bl_int_39_153 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c154
+ bl_int_40_154 bl_int_39_154 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c155
+ bl_int_40_155 bl_int_39_155 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c156
+ bl_int_40_156 bl_int_39_156 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c157
+ bl_int_40_157 bl_int_39_157 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c158
+ bl_int_40_158 bl_int_39_158 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c159
+ bl_int_40_159 bl_int_39_159 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c160
+ bl_int_40_160 bl_int_39_160 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c161
+ bl_int_40_161 bl_int_39_161 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c162
+ bl_int_40_162 bl_int_39_162 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c163
+ bl_int_40_163 bl_int_39_163 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c164
+ bl_int_40_164 bl_int_39_164 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c165
+ bl_int_40_165 bl_int_39_165 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c166
+ bl_int_40_166 bl_int_39_166 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c167
+ bl_int_40_167 bl_int_39_167 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c168
+ bl_int_40_168 bl_int_39_168 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c169
+ bl_int_40_169 bl_int_39_169 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c170
+ bl_int_40_170 bl_int_39_170 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c171
+ bl_int_40_171 bl_int_39_171 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c172
+ bl_int_40_172 bl_int_39_172 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c173
+ bl_int_40_173 bl_int_39_173 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c174
+ bl_int_40_174 bl_int_39_174 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c175
+ bl_int_40_175 bl_int_39_175 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c176
+ bl_int_40_176 bl_int_39_176 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c177
+ bl_int_40_177 bl_int_39_177 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c178
+ bl_int_40_178 bl_int_39_178 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c179
+ bl_int_40_179 bl_int_39_179 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c180
+ bl_int_40_180 bl_int_39_180 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c181
+ bl_int_40_181 bl_int_39_181 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c182
+ bl_int_40_182 bl_int_39_182 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r40_c183
+ bl_int_40_183 bl_int_39_183 wl_0_40 gnd
+ sram_rom_base_one_cell
Xbit_r41_c0
+ bl_int_41_0 bl_int_40_0 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c1
+ bl_int_41_1 bl_int_40_1 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c2
+ bl_int_41_2 bl_int_40_2 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c3
+ bl_int_41_3 bl_int_40_3 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c4
+ bl_int_41_4 bl_int_40_4 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c5
+ bl_int_41_5 bl_int_40_5 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c6
+ bl_int_41_6 bl_int_40_6 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c7
+ bl_int_41_7 bl_int_40_7 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c8
+ bl_int_41_8 bl_int_40_8 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c9
+ bl_int_41_9 bl_int_40_9 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c10
+ bl_int_41_10 bl_int_40_10 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c11
+ bl_int_41_11 bl_int_40_11 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c12
+ bl_int_41_12 bl_int_40_12 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c13
+ bl_int_41_13 bl_int_40_13 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c14
+ bl_int_41_14 bl_int_40_14 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c15
+ bl_int_41_15 bl_int_40_15 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c16
+ bl_int_41_16 bl_int_40_16 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c17
+ bl_int_41_17 bl_int_40_17 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c18
+ bl_int_41_18 bl_int_40_18 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c19
+ bl_int_41_19 bl_int_40_19 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c20
+ bl_int_41_20 bl_int_40_20 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c21
+ bl_int_41_21 bl_int_40_21 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c22
+ bl_int_41_22 bl_int_40_22 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c23
+ bl_int_41_23 bl_int_40_23 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c24
+ bl_int_41_24 bl_int_40_24 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c25
+ bl_int_41_25 bl_int_40_25 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c26
+ bl_int_41_26 bl_int_40_26 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c27
+ bl_int_41_27 bl_int_40_27 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c28
+ bl_int_41_28 bl_int_40_28 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c29
+ bl_int_41_29 bl_int_40_29 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c30
+ bl_int_41_30 bl_int_40_30 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c31
+ bl_int_41_31 bl_int_40_31 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c32
+ bl_int_41_32 bl_int_40_32 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c33
+ bl_int_41_33 bl_int_40_33 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c34
+ bl_int_41_34 bl_int_40_34 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c35
+ bl_int_41_35 bl_int_40_35 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c36
+ bl_int_41_36 bl_int_40_36 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c37
+ bl_int_41_37 bl_int_40_37 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c38
+ bl_int_41_38 bl_int_40_38 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c39
+ bl_int_41_39 bl_int_40_39 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c40
+ bl_int_41_40 bl_int_40_40 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c41
+ bl_int_41_41 bl_int_40_41 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c42
+ bl_int_41_42 bl_int_40_42 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c43
+ bl_int_41_43 bl_int_40_43 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c44
+ bl_int_41_44 bl_int_40_44 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c45
+ bl_int_41_45 bl_int_40_45 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c46
+ bl_int_41_46 bl_int_40_46 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c47
+ bl_int_41_47 bl_int_40_47 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c48
+ bl_int_41_48 bl_int_40_48 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c49
+ bl_int_41_49 bl_int_40_49 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c50
+ bl_int_41_50 bl_int_40_50 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c51
+ bl_int_41_51 bl_int_40_51 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c52
+ bl_int_41_52 bl_int_40_52 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c53
+ bl_int_41_53 bl_int_40_53 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c54
+ bl_int_41_54 bl_int_40_54 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c55
+ bl_int_41_55 bl_int_40_55 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c56
+ bl_int_41_56 bl_int_40_56 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c57
+ bl_int_41_57 bl_int_40_57 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c58
+ bl_int_41_58 bl_int_40_58 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c59
+ bl_int_41_59 bl_int_40_59 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c60
+ bl_int_41_60 bl_int_40_60 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c61
+ bl_int_41_61 bl_int_40_61 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c62
+ bl_int_41_62 bl_int_40_62 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c63
+ bl_int_41_63 bl_int_40_63 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c64
+ bl_int_41_64 bl_int_40_64 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c65
+ bl_int_41_65 bl_int_40_65 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c66
+ bl_int_41_66 bl_int_40_66 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c67
+ bl_int_41_67 bl_int_40_67 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c68
+ bl_int_41_68 bl_int_40_68 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c69
+ bl_int_41_69 bl_int_40_69 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c70
+ bl_int_41_70 bl_int_40_70 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c71
+ bl_int_41_71 bl_int_40_71 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c72
+ bl_int_41_72 bl_int_40_72 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c73
+ bl_int_41_73 bl_int_40_73 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c74
+ bl_int_41_74 bl_int_40_74 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c75
+ bl_int_41_75 bl_int_40_75 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c76
+ bl_int_41_76 bl_int_40_76 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c77
+ bl_int_41_77 bl_int_40_77 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c78
+ bl_int_41_78 bl_int_40_78 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c79
+ bl_int_41_79 bl_int_40_79 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c80
+ bl_int_41_80 bl_int_40_80 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c81
+ bl_int_41_81 bl_int_40_81 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c82
+ bl_int_41_82 bl_int_40_82 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c83
+ bl_int_41_83 bl_int_40_83 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c84
+ bl_int_41_84 bl_int_40_84 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c85
+ bl_int_41_85 bl_int_40_85 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c86
+ bl_int_41_86 bl_int_40_86 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c87
+ bl_int_41_87 bl_int_40_87 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c88
+ bl_int_41_88 bl_int_40_88 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c89
+ bl_int_41_89 bl_int_40_89 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c90
+ bl_int_41_90 bl_int_40_90 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c91
+ bl_int_41_91 bl_int_40_91 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c92
+ bl_int_41_92 bl_int_40_92 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c93
+ bl_int_41_93 bl_int_40_93 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c94
+ bl_int_41_94 bl_int_40_94 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c95
+ bl_int_41_95 bl_int_40_95 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c96
+ bl_int_41_96 bl_int_40_96 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c97
+ bl_int_41_97 bl_int_40_97 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c98
+ bl_int_41_98 bl_int_40_98 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c99
+ bl_int_41_99 bl_int_40_99 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c100
+ bl_int_41_100 bl_int_40_100 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c101
+ bl_int_41_101 bl_int_40_101 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c102
+ bl_int_41_102 bl_int_40_102 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c103
+ bl_int_41_103 bl_int_40_103 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c104
+ bl_int_41_104 bl_int_40_104 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c105
+ bl_int_41_105 bl_int_40_105 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c106
+ bl_int_41_106 bl_int_40_106 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c107
+ bl_int_41_107 bl_int_40_107 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c108
+ bl_int_41_108 bl_int_40_108 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c109
+ bl_int_41_109 bl_int_40_109 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c110
+ bl_int_41_110 bl_int_40_110 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c111
+ bl_int_41_111 bl_int_40_111 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c112
+ bl_int_41_112 bl_int_40_112 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c113
+ bl_int_41_113 bl_int_40_113 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c114
+ bl_int_41_114 bl_int_40_114 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c115
+ bl_int_41_115 bl_int_40_115 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c116
+ bl_int_41_116 bl_int_40_116 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c117
+ bl_int_41_117 bl_int_40_117 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c118
+ bl_int_41_118 bl_int_40_118 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c119
+ bl_int_41_119 bl_int_40_119 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c120
+ bl_int_41_120 bl_int_40_120 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c121
+ bl_int_41_121 bl_int_40_121 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c122
+ bl_int_41_122 bl_int_40_122 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c123
+ bl_int_41_123 bl_int_40_123 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c124
+ bl_int_41_124 bl_int_40_124 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c125
+ bl_int_41_125 bl_int_40_125 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c126
+ bl_int_41_126 bl_int_40_126 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c127
+ bl_int_41_127 bl_int_40_127 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c128
+ bl_int_41_128 bl_int_40_128 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c129
+ bl_int_41_129 bl_int_40_129 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c130
+ bl_int_41_130 bl_int_40_130 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c131
+ bl_int_41_131 bl_int_40_131 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c132
+ bl_int_41_132 bl_int_40_132 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c133
+ bl_int_41_133 bl_int_40_133 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c134
+ bl_int_41_134 bl_int_40_134 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c135
+ bl_int_41_135 bl_int_40_135 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c136
+ bl_int_41_136 bl_int_40_136 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c137
+ bl_int_41_137 bl_int_40_137 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c138
+ bl_int_41_138 bl_int_40_138 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c139
+ bl_int_41_139 bl_int_40_139 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c140
+ bl_int_41_140 bl_int_40_140 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c141
+ bl_int_41_141 bl_int_40_141 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c142
+ bl_int_41_142 bl_int_40_142 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c143
+ bl_int_41_143 bl_int_40_143 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c144
+ bl_int_41_144 bl_int_40_144 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c145
+ bl_int_41_145 bl_int_40_145 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c146
+ bl_int_41_146 bl_int_40_146 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c147
+ bl_int_41_147 bl_int_40_147 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c148
+ bl_int_41_148 bl_int_40_148 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c149
+ bl_int_41_149 bl_int_40_149 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c150
+ bl_int_41_150 bl_int_40_150 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c151
+ bl_int_41_151 bl_int_40_151 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c152
+ bl_int_41_152 bl_int_40_152 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c153
+ bl_int_41_153 bl_int_40_153 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c154
+ bl_int_41_154 bl_int_40_154 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c155
+ bl_int_41_155 bl_int_40_155 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c156
+ bl_int_41_156 bl_int_40_156 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c157
+ bl_int_41_157 bl_int_40_157 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c158
+ bl_int_41_158 bl_int_40_158 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c159
+ bl_int_41_159 bl_int_40_159 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c160
+ bl_int_41_160 bl_int_40_160 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c161
+ bl_int_41_161 bl_int_40_161 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c162
+ bl_int_41_162 bl_int_40_162 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c163
+ bl_int_41_163 bl_int_40_163 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c164
+ bl_int_41_164 bl_int_40_164 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c165
+ bl_int_41_165 bl_int_40_165 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c166
+ bl_int_41_166 bl_int_40_166 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c167
+ bl_int_41_167 bl_int_40_167 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c168
+ bl_int_41_168 bl_int_40_168 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c169
+ bl_int_41_169 bl_int_40_169 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c170
+ bl_int_41_170 bl_int_40_170 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c171
+ bl_int_41_171 bl_int_40_171 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c172
+ bl_int_41_172 bl_int_40_172 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c173
+ bl_int_41_173 bl_int_40_173 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c174
+ bl_int_41_174 bl_int_40_174 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c175
+ bl_int_41_175 bl_int_40_175 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c176
+ bl_int_41_176 bl_int_40_176 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c177
+ bl_int_41_177 bl_int_40_177 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c178
+ bl_int_41_178 bl_int_40_178 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c179
+ bl_int_41_179 bl_int_40_179 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c180
+ bl_int_41_180 bl_int_40_180 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c181
+ bl_int_41_181 bl_int_40_181 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c182
+ bl_int_41_182 bl_int_40_182 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r41_c183
+ bl_int_41_183 bl_int_40_183 wl_0_41 gnd
+ sram_rom_base_one_cell
Xbit_r42_c0
+ bl_int_42_0 bl_int_41_0 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c1
+ bl_int_42_1 bl_int_41_1 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c2
+ bl_int_42_2 bl_int_41_2 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c3
+ bl_int_42_3 bl_int_41_3 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c4
+ bl_int_42_4 bl_int_41_4 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c5
+ bl_int_42_5 bl_int_41_5 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c6
+ bl_int_42_6 bl_int_41_6 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c7
+ bl_int_42_7 bl_int_41_7 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c8
+ bl_int_42_8 bl_int_41_8 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c9
+ bl_int_42_9 bl_int_41_9 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c10
+ bl_int_42_10 bl_int_41_10 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c11
+ bl_int_42_11 bl_int_41_11 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c12
+ bl_int_42_12 bl_int_41_12 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c13
+ bl_int_42_13 bl_int_41_13 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c14
+ bl_int_42_14 bl_int_41_14 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c15
+ bl_int_42_15 bl_int_41_15 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c16
+ bl_int_42_16 bl_int_41_16 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c17
+ bl_int_42_17 bl_int_41_17 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c18
+ bl_int_42_18 bl_int_41_18 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c19
+ bl_int_42_19 bl_int_41_19 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c20
+ bl_int_42_20 bl_int_41_20 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c21
+ bl_int_42_21 bl_int_41_21 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c22
+ bl_int_42_22 bl_int_41_22 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c23
+ bl_int_42_23 bl_int_41_23 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c24
+ bl_int_42_24 bl_int_41_24 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c25
+ bl_int_42_25 bl_int_41_25 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c26
+ bl_int_42_26 bl_int_41_26 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c27
+ bl_int_42_27 bl_int_41_27 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c28
+ bl_int_42_28 bl_int_41_28 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c29
+ bl_int_42_29 bl_int_41_29 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c30
+ bl_int_42_30 bl_int_41_30 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c31
+ bl_int_42_31 bl_int_41_31 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c32
+ bl_int_42_32 bl_int_41_32 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c33
+ bl_int_42_33 bl_int_41_33 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c34
+ bl_int_42_34 bl_int_41_34 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c35
+ bl_int_42_35 bl_int_41_35 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c36
+ bl_int_42_36 bl_int_41_36 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c37
+ bl_int_42_37 bl_int_41_37 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c38
+ bl_int_42_38 bl_int_41_38 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c39
+ bl_int_42_39 bl_int_41_39 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c40
+ bl_int_42_40 bl_int_41_40 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c41
+ bl_int_42_41 bl_int_41_41 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c42
+ bl_int_42_42 bl_int_41_42 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c43
+ bl_int_42_43 bl_int_41_43 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c44
+ bl_int_42_44 bl_int_41_44 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c45
+ bl_int_42_45 bl_int_41_45 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c46
+ bl_int_42_46 bl_int_41_46 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c47
+ bl_int_42_47 bl_int_41_47 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c48
+ bl_int_42_48 bl_int_41_48 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c49
+ bl_int_42_49 bl_int_41_49 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c50
+ bl_int_42_50 bl_int_41_50 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c51
+ bl_int_42_51 bl_int_41_51 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c52
+ bl_int_42_52 bl_int_41_52 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c53
+ bl_int_42_53 bl_int_41_53 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c54
+ bl_int_42_54 bl_int_41_54 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c55
+ bl_int_42_55 bl_int_41_55 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c56
+ bl_int_42_56 bl_int_41_56 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c57
+ bl_int_42_57 bl_int_41_57 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c58
+ bl_int_42_58 bl_int_41_58 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c59
+ bl_int_42_59 bl_int_41_59 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c60
+ bl_int_42_60 bl_int_41_60 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c61
+ bl_int_42_61 bl_int_41_61 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c62
+ bl_int_42_62 bl_int_41_62 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c63
+ bl_int_42_63 bl_int_41_63 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c64
+ bl_int_42_64 bl_int_41_64 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c65
+ bl_int_42_65 bl_int_41_65 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c66
+ bl_int_42_66 bl_int_41_66 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c67
+ bl_int_42_67 bl_int_41_67 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c68
+ bl_int_42_68 bl_int_41_68 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c69
+ bl_int_42_69 bl_int_41_69 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c70
+ bl_int_42_70 bl_int_41_70 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c71
+ bl_int_42_71 bl_int_41_71 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c72
+ bl_int_42_72 bl_int_41_72 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c73
+ bl_int_42_73 bl_int_41_73 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c74
+ bl_int_42_74 bl_int_41_74 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c75
+ bl_int_42_75 bl_int_41_75 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c76
+ bl_int_42_76 bl_int_41_76 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c77
+ bl_int_42_77 bl_int_41_77 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c78
+ bl_int_42_78 bl_int_41_78 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c79
+ bl_int_42_79 bl_int_41_79 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c80
+ bl_int_42_80 bl_int_41_80 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c81
+ bl_int_42_81 bl_int_41_81 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c82
+ bl_int_42_82 bl_int_41_82 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c83
+ bl_int_42_83 bl_int_41_83 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c84
+ bl_int_42_84 bl_int_41_84 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c85
+ bl_int_42_85 bl_int_41_85 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c86
+ bl_int_42_86 bl_int_41_86 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c87
+ bl_int_42_87 bl_int_41_87 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c88
+ bl_int_42_88 bl_int_41_88 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c89
+ bl_int_42_89 bl_int_41_89 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c90
+ bl_int_42_90 bl_int_41_90 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c91
+ bl_int_42_91 bl_int_41_91 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c92
+ bl_int_42_92 bl_int_41_92 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c93
+ bl_int_42_93 bl_int_41_93 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c94
+ bl_int_42_94 bl_int_41_94 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c95
+ bl_int_42_95 bl_int_41_95 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c96
+ bl_int_42_96 bl_int_41_96 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c97
+ bl_int_42_97 bl_int_41_97 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c98
+ bl_int_42_98 bl_int_41_98 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c99
+ bl_int_42_99 bl_int_41_99 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c100
+ bl_int_42_100 bl_int_41_100 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c101
+ bl_int_42_101 bl_int_41_101 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c102
+ bl_int_42_102 bl_int_41_102 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c103
+ bl_int_42_103 bl_int_41_103 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c104
+ bl_int_42_104 bl_int_41_104 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c105
+ bl_int_42_105 bl_int_41_105 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c106
+ bl_int_42_106 bl_int_41_106 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c107
+ bl_int_42_107 bl_int_41_107 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c108
+ bl_int_42_108 bl_int_41_108 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c109
+ bl_int_42_109 bl_int_41_109 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c110
+ bl_int_42_110 bl_int_41_110 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c111
+ bl_int_42_111 bl_int_41_111 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c112
+ bl_int_42_112 bl_int_41_112 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c113
+ bl_int_42_113 bl_int_41_113 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c114
+ bl_int_42_114 bl_int_41_114 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c115
+ bl_int_42_115 bl_int_41_115 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c116
+ bl_int_42_116 bl_int_41_116 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c117
+ bl_int_42_117 bl_int_41_117 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c118
+ bl_int_42_118 bl_int_41_118 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c119
+ bl_int_42_119 bl_int_41_119 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c120
+ bl_int_42_120 bl_int_41_120 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c121
+ bl_int_42_121 bl_int_41_121 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c122
+ bl_int_42_122 bl_int_41_122 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c123
+ bl_int_42_123 bl_int_41_123 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c124
+ bl_int_42_124 bl_int_41_124 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c125
+ bl_int_42_125 bl_int_41_125 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c126
+ bl_int_42_126 bl_int_41_126 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c127
+ bl_int_42_127 bl_int_41_127 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c128
+ bl_int_42_128 bl_int_41_128 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c129
+ bl_int_42_129 bl_int_41_129 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c130
+ bl_int_42_130 bl_int_41_130 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c131
+ bl_int_42_131 bl_int_41_131 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c132
+ bl_int_42_132 bl_int_41_132 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c133
+ bl_int_42_133 bl_int_41_133 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c134
+ bl_int_42_134 bl_int_41_134 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c135
+ bl_int_42_135 bl_int_41_135 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c136
+ bl_int_42_136 bl_int_41_136 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c137
+ bl_int_42_137 bl_int_41_137 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c138
+ bl_int_42_138 bl_int_41_138 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c139
+ bl_int_42_139 bl_int_41_139 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c140
+ bl_int_42_140 bl_int_41_140 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c141
+ bl_int_42_141 bl_int_41_141 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c142
+ bl_int_42_142 bl_int_41_142 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c143
+ bl_int_42_143 bl_int_41_143 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c144
+ bl_int_42_144 bl_int_41_144 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c145
+ bl_int_42_145 bl_int_41_145 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c146
+ bl_int_42_146 bl_int_41_146 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c147
+ bl_int_42_147 bl_int_41_147 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c148
+ bl_int_42_148 bl_int_41_148 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c149
+ bl_int_42_149 bl_int_41_149 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c150
+ bl_int_42_150 bl_int_41_150 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c151
+ bl_int_42_151 bl_int_41_151 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c152
+ bl_int_42_152 bl_int_41_152 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c153
+ bl_int_42_153 bl_int_41_153 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c154
+ bl_int_42_154 bl_int_41_154 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c155
+ bl_int_42_155 bl_int_41_155 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c156
+ bl_int_42_156 bl_int_41_156 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c157
+ bl_int_42_157 bl_int_41_157 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c158
+ bl_int_42_158 bl_int_41_158 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c159
+ bl_int_42_159 bl_int_41_159 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c160
+ bl_int_42_160 bl_int_41_160 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c161
+ bl_int_42_161 bl_int_41_161 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c162
+ bl_int_42_162 bl_int_41_162 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c163
+ bl_int_42_163 bl_int_41_163 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c164
+ bl_int_42_164 bl_int_41_164 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c165
+ bl_int_42_165 bl_int_41_165 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c166
+ bl_int_42_166 bl_int_41_166 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c167
+ bl_int_42_167 bl_int_41_167 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c168
+ bl_int_42_168 bl_int_41_168 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c169
+ bl_int_42_169 bl_int_41_169 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c170
+ bl_int_42_170 bl_int_41_170 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c171
+ bl_int_42_171 bl_int_41_171 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c172
+ bl_int_42_172 bl_int_41_172 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c173
+ bl_int_42_173 bl_int_41_173 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c174
+ bl_int_42_174 bl_int_41_174 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c175
+ bl_int_42_175 bl_int_41_175 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c176
+ bl_int_42_176 bl_int_41_176 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c177
+ bl_int_42_177 bl_int_41_177 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c178
+ bl_int_42_178 bl_int_41_178 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c179
+ bl_int_42_179 bl_int_41_179 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c180
+ bl_int_42_180 bl_int_41_180 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c181
+ bl_int_42_181 bl_int_41_181 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c182
+ bl_int_42_182 bl_int_41_182 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r42_c183
+ bl_int_42_183 bl_int_41_183 wl_0_42 gnd
+ sram_rom_base_one_cell
Xbit_r43_c0
+ bl_int_43_0 bl_int_42_0 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c1
+ bl_int_43_1 bl_int_42_1 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c2
+ bl_int_43_2 bl_int_42_2 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c3
+ bl_int_42_3 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c4
+ bl_int_42_4 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c5
+ bl_int_42_5 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c6
+ bl_int_42_6 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c7
+ bl_int_42_7 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c8
+ bl_int_42_8 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c9
+ bl_int_42_9 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c10
+ bl_int_42_10 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c11
+ bl_int_42_11 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c12
+ bl_int_42_12 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c13
+ bl_int_42_13 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c14
+ bl_int_42_14 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c15
+ bl_int_42_15 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c16
+ bl_int_42_16 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c17
+ bl_int_42_17 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c18
+ bl_int_42_18 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c19
+ bl_int_43_19 bl_int_42_19 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c20
+ bl_int_43_20 bl_int_42_20 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c21
+ bl_int_43_21 bl_int_42_21 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c22
+ bl_int_43_22 bl_int_42_22 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c23
+ bl_int_43_23 bl_int_42_23 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c24
+ bl_int_43_24 bl_int_42_24 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c25
+ bl_int_43_25 bl_int_42_25 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c26
+ bl_int_42_26 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c27
+ bl_int_42_27 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c28
+ bl_int_42_28 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c29
+ bl_int_42_29 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c30
+ bl_int_42_30 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c31
+ bl_int_42_31 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c32
+ bl_int_42_32 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c33
+ bl_int_42_33 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c34
+ bl_int_42_34 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c35
+ bl_int_42_35 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c36
+ bl_int_42_36 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c37
+ bl_int_42_37 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c38
+ bl_int_42_38 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c39
+ bl_int_42_39 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c40
+ bl_int_42_40 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c41
+ bl_int_42_41 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c42
+ bl_int_43_42 bl_int_42_42 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c43
+ bl_int_43_43 bl_int_42_43 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c44
+ bl_int_43_44 bl_int_42_44 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c45
+ bl_int_43_45 bl_int_42_45 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c46
+ bl_int_43_46 bl_int_42_46 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c47
+ bl_int_43_47 bl_int_42_47 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c48
+ bl_int_43_48 bl_int_42_48 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c49
+ bl_int_42_49 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c50
+ bl_int_42_50 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c51
+ bl_int_42_51 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c52
+ bl_int_42_52 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c53
+ bl_int_42_53 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c54
+ bl_int_42_54 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c55
+ bl_int_42_55 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c56
+ bl_int_42_56 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c57
+ bl_int_42_57 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c58
+ bl_int_42_58 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c59
+ bl_int_42_59 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c60
+ bl_int_42_60 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c61
+ bl_int_42_61 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c62
+ bl_int_42_62 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c63
+ bl_int_42_63 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c64
+ bl_int_42_64 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c65
+ bl_int_43_65 bl_int_42_65 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c66
+ bl_int_43_66 bl_int_42_66 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c67
+ bl_int_43_67 bl_int_42_67 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c68
+ bl_int_43_68 bl_int_42_68 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c69
+ bl_int_43_69 bl_int_42_69 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c70
+ bl_int_43_70 bl_int_42_70 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c71
+ bl_int_43_71 bl_int_42_71 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c72
+ bl_int_42_72 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c73
+ bl_int_42_73 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c74
+ bl_int_42_74 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c75
+ bl_int_42_75 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c76
+ bl_int_42_76 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c77
+ bl_int_42_77 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c78
+ bl_int_42_78 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c79
+ bl_int_42_79 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c80
+ bl_int_42_80 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c81
+ bl_int_42_81 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c82
+ bl_int_42_82 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c83
+ bl_int_42_83 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c84
+ bl_int_42_84 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c85
+ bl_int_42_85 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c86
+ bl_int_42_86 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c87
+ bl_int_42_87 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c88
+ bl_int_43_88 bl_int_42_88 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c89
+ bl_int_43_89 bl_int_42_89 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c90
+ bl_int_43_90 bl_int_42_90 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c91
+ bl_int_43_91 bl_int_42_91 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c92
+ bl_int_43_92 bl_int_42_92 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c93
+ bl_int_43_93 bl_int_42_93 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c94
+ bl_int_43_94 bl_int_42_94 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c95
+ bl_int_42_95 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c96
+ bl_int_42_96 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c97
+ bl_int_42_97 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c98
+ bl_int_42_98 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c99
+ bl_int_42_99 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c100
+ bl_int_42_100 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c101
+ bl_int_42_101 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c102
+ bl_int_42_102 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c103
+ bl_int_42_103 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c104
+ bl_int_42_104 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c105
+ bl_int_42_105 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c106
+ bl_int_42_106 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c107
+ bl_int_42_107 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c108
+ bl_int_42_108 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c109
+ bl_int_42_109 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c110
+ bl_int_42_110 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c111
+ bl_int_43_111 bl_int_42_111 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c112
+ bl_int_43_112 bl_int_42_112 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c113
+ bl_int_43_113 bl_int_42_113 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c114
+ bl_int_43_114 bl_int_42_114 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c115
+ bl_int_43_115 bl_int_42_115 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c116
+ bl_int_43_116 bl_int_42_116 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c117
+ bl_int_43_117 bl_int_42_117 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c118
+ bl_int_42_118 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c119
+ bl_int_42_119 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c120
+ bl_int_42_120 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c121
+ bl_int_42_121 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c122
+ bl_int_42_122 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c123
+ bl_int_42_123 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c124
+ bl_int_42_124 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c125
+ bl_int_42_125 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c126
+ bl_int_42_126 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c127
+ bl_int_42_127 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c128
+ bl_int_42_128 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c129
+ bl_int_42_129 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c130
+ bl_int_42_130 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c131
+ bl_int_42_131 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c132
+ bl_int_42_132 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c133
+ bl_int_42_133 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c134
+ bl_int_43_134 bl_int_42_134 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c135
+ bl_int_43_135 bl_int_42_135 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c136
+ bl_int_43_136 bl_int_42_136 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c137
+ bl_int_43_137 bl_int_42_137 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c138
+ bl_int_43_138 bl_int_42_138 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c139
+ bl_int_43_139 bl_int_42_139 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c140
+ bl_int_43_140 bl_int_42_140 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c141
+ bl_int_42_141 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c142
+ bl_int_42_142 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c143
+ bl_int_42_143 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c144
+ bl_int_42_144 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c145
+ bl_int_42_145 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c146
+ bl_int_42_146 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c147
+ bl_int_42_147 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c148
+ bl_int_42_148 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c149
+ bl_int_42_149 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c150
+ bl_int_42_150 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c151
+ bl_int_42_151 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c152
+ bl_int_42_152 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c153
+ bl_int_42_153 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c154
+ bl_int_42_154 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c155
+ bl_int_42_155 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c156
+ bl_int_42_156 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c157
+ bl_int_43_157 bl_int_42_157 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c158
+ bl_int_43_158 bl_int_42_158 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c159
+ bl_int_43_159 bl_int_42_159 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c160
+ bl_int_43_160 bl_int_42_160 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c161
+ bl_int_43_161 bl_int_42_161 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c162
+ bl_int_43_162 bl_int_42_162 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c163
+ bl_int_43_163 bl_int_42_163 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c164
+ bl_int_42_164 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c165
+ bl_int_42_165 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c166
+ bl_int_42_166 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c167
+ bl_int_42_167 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c168
+ bl_int_42_168 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c169
+ bl_int_42_169 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c170
+ bl_int_42_170 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c171
+ bl_int_42_171 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c172
+ bl_int_42_172 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c173
+ bl_int_42_173 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c174
+ bl_int_42_174 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c175
+ bl_int_42_175 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c176
+ bl_int_42_176 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c177
+ bl_int_42_177 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c178
+ bl_int_42_178 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c179
+ bl_int_42_179 wl_0_43 gnd
+ sram_rom_base_zero_cell
Xbit_r43_c180
+ bl_int_43_180 bl_int_42_180 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c181
+ bl_int_43_181 bl_int_42_181 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c182
+ bl_int_43_182 bl_int_42_182 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r43_c183
+ bl_int_43_183 bl_int_42_183 wl_0_43 gnd
+ sram_rom_base_one_cell
Xbit_r44_c0
+ bl_int_44_0 bl_int_43_0 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c1
+ bl_int_44_1 bl_int_43_1 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c2
+ bl_int_44_2 bl_int_43_2 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c3
+ bl_int_44_3 bl_int_42_3 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c4
+ bl_int_44_4 bl_int_42_4 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c5
+ bl_int_44_5 bl_int_42_5 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c6
+ bl_int_44_6 bl_int_42_6 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c7
+ bl_int_44_7 bl_int_42_7 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c8
+ bl_int_44_8 bl_int_42_8 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c9
+ bl_int_44_9 bl_int_42_9 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c10
+ bl_int_44_10 bl_int_42_10 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c11
+ bl_int_44_11 bl_int_42_11 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c12
+ bl_int_44_12 bl_int_42_12 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c13
+ bl_int_44_13 bl_int_42_13 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c14
+ bl_int_44_14 bl_int_42_14 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c15
+ bl_int_44_15 bl_int_42_15 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c16
+ bl_int_44_16 bl_int_42_16 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c17
+ bl_int_44_17 bl_int_42_17 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c18
+ bl_int_44_18 bl_int_42_18 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c19
+ bl_int_44_19 bl_int_43_19 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c20
+ bl_int_44_20 bl_int_43_20 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c21
+ bl_int_44_21 bl_int_43_21 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c22
+ bl_int_44_22 bl_int_43_22 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c23
+ bl_int_44_23 bl_int_43_23 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c24
+ bl_int_44_24 bl_int_43_24 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c25
+ bl_int_44_25 bl_int_43_25 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c26
+ bl_int_44_26 bl_int_42_26 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c27
+ bl_int_44_27 bl_int_42_27 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c28
+ bl_int_44_28 bl_int_42_28 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c29
+ bl_int_44_29 bl_int_42_29 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c30
+ bl_int_44_30 bl_int_42_30 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c31
+ bl_int_44_31 bl_int_42_31 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c32
+ bl_int_44_32 bl_int_42_32 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c33
+ bl_int_44_33 bl_int_42_33 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c34
+ bl_int_44_34 bl_int_42_34 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c35
+ bl_int_44_35 bl_int_42_35 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c36
+ bl_int_44_36 bl_int_42_36 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c37
+ bl_int_44_37 bl_int_42_37 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c38
+ bl_int_44_38 bl_int_42_38 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c39
+ bl_int_44_39 bl_int_42_39 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c40
+ bl_int_44_40 bl_int_42_40 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c41
+ bl_int_44_41 bl_int_42_41 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c42
+ bl_int_44_42 bl_int_43_42 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c43
+ bl_int_44_43 bl_int_43_43 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c44
+ bl_int_44_44 bl_int_43_44 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c45
+ bl_int_44_45 bl_int_43_45 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c46
+ bl_int_44_46 bl_int_43_46 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c47
+ bl_int_44_47 bl_int_43_47 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c48
+ bl_int_44_48 bl_int_43_48 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c49
+ bl_int_44_49 bl_int_42_49 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c50
+ bl_int_44_50 bl_int_42_50 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c51
+ bl_int_44_51 bl_int_42_51 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c52
+ bl_int_44_52 bl_int_42_52 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c53
+ bl_int_44_53 bl_int_42_53 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c54
+ bl_int_44_54 bl_int_42_54 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c55
+ bl_int_44_55 bl_int_42_55 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c56
+ bl_int_44_56 bl_int_42_56 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c57
+ bl_int_44_57 bl_int_42_57 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c58
+ bl_int_44_58 bl_int_42_58 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c59
+ bl_int_44_59 bl_int_42_59 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c60
+ bl_int_44_60 bl_int_42_60 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c61
+ bl_int_44_61 bl_int_42_61 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c62
+ bl_int_44_62 bl_int_42_62 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c63
+ bl_int_44_63 bl_int_42_63 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c64
+ bl_int_44_64 bl_int_42_64 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c65
+ bl_int_44_65 bl_int_43_65 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c66
+ bl_int_44_66 bl_int_43_66 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c67
+ bl_int_44_67 bl_int_43_67 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c68
+ bl_int_44_68 bl_int_43_68 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c69
+ bl_int_44_69 bl_int_43_69 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c70
+ bl_int_44_70 bl_int_43_70 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c71
+ bl_int_44_71 bl_int_43_71 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c72
+ bl_int_44_72 bl_int_42_72 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c73
+ bl_int_44_73 bl_int_42_73 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c74
+ bl_int_44_74 bl_int_42_74 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c75
+ bl_int_44_75 bl_int_42_75 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c76
+ bl_int_44_76 bl_int_42_76 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c77
+ bl_int_44_77 bl_int_42_77 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c78
+ bl_int_44_78 bl_int_42_78 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c79
+ bl_int_44_79 bl_int_42_79 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c80
+ bl_int_44_80 bl_int_42_80 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c81
+ bl_int_44_81 bl_int_42_81 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c82
+ bl_int_44_82 bl_int_42_82 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c83
+ bl_int_44_83 bl_int_42_83 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c84
+ bl_int_44_84 bl_int_42_84 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c85
+ bl_int_44_85 bl_int_42_85 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c86
+ bl_int_44_86 bl_int_42_86 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c87
+ bl_int_44_87 bl_int_42_87 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c88
+ bl_int_44_88 bl_int_43_88 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c89
+ bl_int_44_89 bl_int_43_89 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c90
+ bl_int_44_90 bl_int_43_90 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c91
+ bl_int_44_91 bl_int_43_91 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c92
+ bl_int_44_92 bl_int_43_92 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c93
+ bl_int_44_93 bl_int_43_93 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c94
+ bl_int_44_94 bl_int_43_94 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c95
+ bl_int_44_95 bl_int_42_95 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c96
+ bl_int_44_96 bl_int_42_96 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c97
+ bl_int_44_97 bl_int_42_97 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c98
+ bl_int_44_98 bl_int_42_98 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c99
+ bl_int_44_99 bl_int_42_99 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c100
+ bl_int_44_100 bl_int_42_100 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c101
+ bl_int_44_101 bl_int_42_101 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c102
+ bl_int_44_102 bl_int_42_102 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c103
+ bl_int_44_103 bl_int_42_103 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c104
+ bl_int_44_104 bl_int_42_104 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c105
+ bl_int_44_105 bl_int_42_105 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c106
+ bl_int_44_106 bl_int_42_106 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c107
+ bl_int_44_107 bl_int_42_107 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c108
+ bl_int_44_108 bl_int_42_108 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c109
+ bl_int_44_109 bl_int_42_109 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c110
+ bl_int_44_110 bl_int_42_110 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c111
+ bl_int_44_111 bl_int_43_111 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c112
+ bl_int_44_112 bl_int_43_112 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c113
+ bl_int_44_113 bl_int_43_113 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c114
+ bl_int_44_114 bl_int_43_114 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c115
+ bl_int_44_115 bl_int_43_115 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c116
+ bl_int_44_116 bl_int_43_116 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c117
+ bl_int_44_117 bl_int_43_117 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c118
+ bl_int_44_118 bl_int_42_118 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c119
+ bl_int_44_119 bl_int_42_119 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c120
+ bl_int_44_120 bl_int_42_120 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c121
+ bl_int_44_121 bl_int_42_121 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c122
+ bl_int_44_122 bl_int_42_122 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c123
+ bl_int_44_123 bl_int_42_123 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c124
+ bl_int_44_124 bl_int_42_124 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c125
+ bl_int_44_125 bl_int_42_125 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c126
+ bl_int_44_126 bl_int_42_126 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c127
+ bl_int_44_127 bl_int_42_127 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c128
+ bl_int_44_128 bl_int_42_128 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c129
+ bl_int_44_129 bl_int_42_129 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c130
+ bl_int_44_130 bl_int_42_130 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c131
+ bl_int_44_131 bl_int_42_131 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c132
+ bl_int_44_132 bl_int_42_132 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c133
+ bl_int_44_133 bl_int_42_133 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c134
+ bl_int_44_134 bl_int_43_134 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c135
+ bl_int_44_135 bl_int_43_135 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c136
+ bl_int_44_136 bl_int_43_136 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c137
+ bl_int_44_137 bl_int_43_137 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c138
+ bl_int_44_138 bl_int_43_138 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c139
+ bl_int_44_139 bl_int_43_139 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c140
+ bl_int_44_140 bl_int_43_140 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c141
+ bl_int_44_141 bl_int_42_141 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c142
+ bl_int_44_142 bl_int_42_142 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c143
+ bl_int_44_143 bl_int_42_143 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c144
+ bl_int_44_144 bl_int_42_144 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c145
+ bl_int_44_145 bl_int_42_145 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c146
+ bl_int_44_146 bl_int_42_146 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c147
+ bl_int_44_147 bl_int_42_147 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c148
+ bl_int_44_148 bl_int_42_148 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c149
+ bl_int_44_149 bl_int_42_149 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c150
+ bl_int_44_150 bl_int_42_150 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c151
+ bl_int_44_151 bl_int_42_151 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c152
+ bl_int_44_152 bl_int_42_152 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c153
+ bl_int_44_153 bl_int_42_153 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c154
+ bl_int_44_154 bl_int_42_154 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c155
+ bl_int_44_155 bl_int_42_155 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c156
+ bl_int_44_156 bl_int_42_156 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c157
+ bl_int_44_157 bl_int_43_157 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c158
+ bl_int_44_158 bl_int_43_158 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c159
+ bl_int_44_159 bl_int_43_159 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c160
+ bl_int_44_160 bl_int_43_160 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c161
+ bl_int_44_161 bl_int_43_161 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c162
+ bl_int_44_162 bl_int_43_162 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c163
+ bl_int_44_163 bl_int_43_163 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c164
+ bl_int_44_164 bl_int_42_164 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c165
+ bl_int_44_165 bl_int_42_165 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c166
+ bl_int_44_166 bl_int_42_166 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c167
+ bl_int_44_167 bl_int_42_167 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c168
+ bl_int_44_168 bl_int_42_168 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c169
+ bl_int_44_169 bl_int_42_169 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c170
+ bl_int_44_170 bl_int_42_170 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c171
+ bl_int_44_171 bl_int_42_171 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c172
+ bl_int_44_172 bl_int_42_172 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c173
+ bl_int_44_173 bl_int_42_173 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c174
+ bl_int_44_174 bl_int_42_174 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c175
+ bl_int_44_175 bl_int_42_175 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c176
+ bl_int_44_176 bl_int_42_176 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c177
+ bl_int_44_177 bl_int_42_177 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c178
+ bl_int_44_178 bl_int_42_178 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c179
+ bl_int_44_179 bl_int_42_179 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c180
+ bl_int_44_180 bl_int_43_180 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c181
+ bl_int_44_181 bl_int_43_181 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c182
+ bl_int_44_182 bl_int_43_182 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r44_c183
+ bl_int_44_183 bl_int_43_183 wl_0_44 gnd
+ sram_rom_base_one_cell
Xbit_r45_c0
+ bl_int_45_0 bl_int_44_0 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c1
+ bl_int_45_1 bl_int_44_1 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c2
+ bl_int_45_2 bl_int_44_2 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c3
+ bl_int_45_3 bl_int_44_3 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c4
+ bl_int_45_4 bl_int_44_4 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c5
+ bl_int_45_5 bl_int_44_5 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c6
+ bl_int_45_6 bl_int_44_6 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c7
+ bl_int_45_7 bl_int_44_7 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c8
+ bl_int_45_8 bl_int_44_8 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c9
+ bl_int_45_9 bl_int_44_9 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c10
+ bl_int_45_10 bl_int_44_10 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c11
+ bl_int_45_11 bl_int_44_11 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c12
+ bl_int_45_12 bl_int_44_12 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c13
+ bl_int_45_13 bl_int_44_13 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c14
+ bl_int_45_14 bl_int_44_14 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c15
+ bl_int_45_15 bl_int_44_15 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c16
+ bl_int_45_16 bl_int_44_16 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c17
+ bl_int_45_17 bl_int_44_17 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c18
+ bl_int_45_18 bl_int_44_18 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c19
+ bl_int_45_19 bl_int_44_19 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c20
+ bl_int_45_20 bl_int_44_20 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c21
+ bl_int_45_21 bl_int_44_21 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c22
+ bl_int_45_22 bl_int_44_22 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c23
+ bl_int_45_23 bl_int_44_23 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c24
+ bl_int_45_24 bl_int_44_24 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c25
+ bl_int_45_25 bl_int_44_25 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c26
+ bl_int_45_26 bl_int_44_26 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c27
+ bl_int_45_27 bl_int_44_27 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c28
+ bl_int_45_28 bl_int_44_28 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c29
+ bl_int_45_29 bl_int_44_29 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c30
+ bl_int_45_30 bl_int_44_30 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c31
+ bl_int_45_31 bl_int_44_31 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c32
+ bl_int_45_32 bl_int_44_32 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c33
+ bl_int_45_33 bl_int_44_33 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c34
+ bl_int_45_34 bl_int_44_34 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c35
+ bl_int_45_35 bl_int_44_35 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c36
+ bl_int_45_36 bl_int_44_36 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c37
+ bl_int_45_37 bl_int_44_37 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c38
+ bl_int_45_38 bl_int_44_38 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c39
+ bl_int_45_39 bl_int_44_39 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c40
+ bl_int_45_40 bl_int_44_40 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c41
+ bl_int_45_41 bl_int_44_41 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c42
+ bl_int_45_42 bl_int_44_42 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c43
+ bl_int_45_43 bl_int_44_43 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c44
+ bl_int_45_44 bl_int_44_44 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c45
+ bl_int_45_45 bl_int_44_45 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c46
+ bl_int_45_46 bl_int_44_46 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c47
+ bl_int_45_47 bl_int_44_47 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c48
+ bl_int_45_48 bl_int_44_48 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c49
+ bl_int_45_49 bl_int_44_49 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c50
+ bl_int_45_50 bl_int_44_50 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c51
+ bl_int_45_51 bl_int_44_51 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c52
+ bl_int_45_52 bl_int_44_52 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c53
+ bl_int_45_53 bl_int_44_53 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c54
+ bl_int_45_54 bl_int_44_54 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c55
+ bl_int_45_55 bl_int_44_55 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c56
+ bl_int_45_56 bl_int_44_56 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c57
+ bl_int_45_57 bl_int_44_57 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c58
+ bl_int_45_58 bl_int_44_58 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c59
+ bl_int_45_59 bl_int_44_59 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c60
+ bl_int_45_60 bl_int_44_60 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c61
+ bl_int_45_61 bl_int_44_61 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c62
+ bl_int_45_62 bl_int_44_62 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c63
+ bl_int_45_63 bl_int_44_63 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c64
+ bl_int_45_64 bl_int_44_64 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c65
+ bl_int_45_65 bl_int_44_65 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c66
+ bl_int_45_66 bl_int_44_66 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c67
+ bl_int_45_67 bl_int_44_67 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c68
+ bl_int_45_68 bl_int_44_68 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c69
+ bl_int_45_69 bl_int_44_69 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c70
+ bl_int_45_70 bl_int_44_70 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c71
+ bl_int_45_71 bl_int_44_71 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c72
+ bl_int_45_72 bl_int_44_72 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c73
+ bl_int_45_73 bl_int_44_73 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c74
+ bl_int_45_74 bl_int_44_74 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c75
+ bl_int_45_75 bl_int_44_75 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c76
+ bl_int_45_76 bl_int_44_76 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c77
+ bl_int_45_77 bl_int_44_77 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c78
+ bl_int_45_78 bl_int_44_78 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c79
+ bl_int_45_79 bl_int_44_79 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c80
+ bl_int_45_80 bl_int_44_80 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c81
+ bl_int_45_81 bl_int_44_81 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c82
+ bl_int_45_82 bl_int_44_82 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c83
+ bl_int_45_83 bl_int_44_83 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c84
+ bl_int_45_84 bl_int_44_84 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c85
+ bl_int_45_85 bl_int_44_85 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c86
+ bl_int_45_86 bl_int_44_86 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c87
+ bl_int_45_87 bl_int_44_87 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c88
+ bl_int_45_88 bl_int_44_88 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c89
+ bl_int_45_89 bl_int_44_89 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c90
+ bl_int_45_90 bl_int_44_90 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c91
+ bl_int_45_91 bl_int_44_91 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c92
+ bl_int_45_92 bl_int_44_92 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c93
+ bl_int_45_93 bl_int_44_93 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c94
+ bl_int_45_94 bl_int_44_94 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c95
+ bl_int_45_95 bl_int_44_95 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c96
+ bl_int_45_96 bl_int_44_96 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c97
+ bl_int_45_97 bl_int_44_97 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c98
+ bl_int_45_98 bl_int_44_98 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c99
+ bl_int_45_99 bl_int_44_99 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c100
+ bl_int_45_100 bl_int_44_100 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c101
+ bl_int_45_101 bl_int_44_101 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c102
+ bl_int_45_102 bl_int_44_102 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c103
+ bl_int_45_103 bl_int_44_103 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c104
+ bl_int_45_104 bl_int_44_104 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c105
+ bl_int_45_105 bl_int_44_105 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c106
+ bl_int_45_106 bl_int_44_106 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c107
+ bl_int_45_107 bl_int_44_107 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c108
+ bl_int_45_108 bl_int_44_108 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c109
+ bl_int_45_109 bl_int_44_109 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c110
+ bl_int_45_110 bl_int_44_110 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c111
+ bl_int_45_111 bl_int_44_111 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c112
+ bl_int_45_112 bl_int_44_112 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c113
+ bl_int_45_113 bl_int_44_113 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c114
+ bl_int_45_114 bl_int_44_114 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c115
+ bl_int_45_115 bl_int_44_115 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c116
+ bl_int_45_116 bl_int_44_116 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c117
+ bl_int_45_117 bl_int_44_117 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c118
+ bl_int_45_118 bl_int_44_118 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c119
+ bl_int_45_119 bl_int_44_119 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c120
+ bl_int_45_120 bl_int_44_120 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c121
+ bl_int_45_121 bl_int_44_121 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c122
+ bl_int_45_122 bl_int_44_122 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c123
+ bl_int_45_123 bl_int_44_123 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c124
+ bl_int_45_124 bl_int_44_124 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c125
+ bl_int_45_125 bl_int_44_125 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c126
+ bl_int_45_126 bl_int_44_126 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c127
+ bl_int_45_127 bl_int_44_127 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c128
+ bl_int_45_128 bl_int_44_128 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c129
+ bl_int_45_129 bl_int_44_129 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c130
+ bl_int_45_130 bl_int_44_130 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c131
+ bl_int_45_131 bl_int_44_131 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c132
+ bl_int_45_132 bl_int_44_132 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c133
+ bl_int_45_133 bl_int_44_133 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c134
+ bl_int_45_134 bl_int_44_134 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c135
+ bl_int_45_135 bl_int_44_135 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c136
+ bl_int_45_136 bl_int_44_136 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c137
+ bl_int_45_137 bl_int_44_137 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c138
+ bl_int_45_138 bl_int_44_138 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c139
+ bl_int_45_139 bl_int_44_139 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c140
+ bl_int_45_140 bl_int_44_140 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c141
+ bl_int_45_141 bl_int_44_141 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c142
+ bl_int_45_142 bl_int_44_142 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c143
+ bl_int_45_143 bl_int_44_143 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c144
+ bl_int_45_144 bl_int_44_144 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c145
+ bl_int_45_145 bl_int_44_145 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c146
+ bl_int_45_146 bl_int_44_146 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c147
+ bl_int_45_147 bl_int_44_147 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c148
+ bl_int_45_148 bl_int_44_148 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c149
+ bl_int_45_149 bl_int_44_149 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c150
+ bl_int_45_150 bl_int_44_150 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c151
+ bl_int_45_151 bl_int_44_151 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c152
+ bl_int_45_152 bl_int_44_152 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c153
+ bl_int_45_153 bl_int_44_153 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c154
+ bl_int_45_154 bl_int_44_154 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c155
+ bl_int_45_155 bl_int_44_155 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c156
+ bl_int_45_156 bl_int_44_156 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c157
+ bl_int_45_157 bl_int_44_157 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c158
+ bl_int_45_158 bl_int_44_158 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c159
+ bl_int_45_159 bl_int_44_159 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c160
+ bl_int_45_160 bl_int_44_160 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c161
+ bl_int_45_161 bl_int_44_161 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c162
+ bl_int_45_162 bl_int_44_162 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c163
+ bl_int_45_163 bl_int_44_163 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c164
+ bl_int_45_164 bl_int_44_164 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c165
+ bl_int_45_165 bl_int_44_165 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c166
+ bl_int_45_166 bl_int_44_166 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c167
+ bl_int_45_167 bl_int_44_167 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c168
+ bl_int_45_168 bl_int_44_168 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c169
+ bl_int_45_169 bl_int_44_169 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c170
+ bl_int_45_170 bl_int_44_170 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c171
+ bl_int_45_171 bl_int_44_171 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c172
+ bl_int_45_172 bl_int_44_172 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c173
+ bl_int_45_173 bl_int_44_173 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c174
+ bl_int_45_174 bl_int_44_174 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c175
+ bl_int_45_175 bl_int_44_175 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c176
+ bl_int_45_176 bl_int_44_176 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c177
+ bl_int_45_177 bl_int_44_177 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c178
+ bl_int_45_178 bl_int_44_178 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c179
+ bl_int_45_179 bl_int_44_179 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c180
+ bl_int_45_180 bl_int_44_180 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c181
+ bl_int_45_181 bl_int_44_181 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c182
+ bl_int_45_182 bl_int_44_182 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r45_c183
+ bl_int_45_183 bl_int_44_183 wl_0_45 gnd
+ sram_rom_base_one_cell
Xbit_r46_c0
+ bl_int_46_0 bl_int_45_0 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c1
+ bl_int_46_1 bl_int_45_1 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c2
+ bl_int_46_2 bl_int_45_2 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c3
+ bl_int_46_3 bl_int_45_3 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c4
+ bl_int_46_4 bl_int_45_4 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c5
+ bl_int_46_5 bl_int_45_5 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c6
+ bl_int_46_6 bl_int_45_6 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c7
+ bl_int_46_7 bl_int_45_7 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c8
+ bl_int_46_8 bl_int_45_8 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c9
+ bl_int_46_9 bl_int_45_9 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c10
+ bl_int_46_10 bl_int_45_10 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c11
+ bl_int_46_11 bl_int_45_11 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c12
+ bl_int_46_12 bl_int_45_12 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c13
+ bl_int_46_13 bl_int_45_13 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c14
+ bl_int_46_14 bl_int_45_14 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c15
+ bl_int_46_15 bl_int_45_15 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c16
+ bl_int_46_16 bl_int_45_16 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c17
+ bl_int_46_17 bl_int_45_17 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c18
+ bl_int_46_18 bl_int_45_18 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c19
+ bl_int_46_19 bl_int_45_19 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c20
+ bl_int_46_20 bl_int_45_20 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c21
+ bl_int_46_21 bl_int_45_21 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c22
+ bl_int_46_22 bl_int_45_22 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c23
+ bl_int_46_23 bl_int_45_23 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c24
+ bl_int_46_24 bl_int_45_24 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c25
+ bl_int_46_25 bl_int_45_25 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c26
+ bl_int_46_26 bl_int_45_26 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c27
+ bl_int_46_27 bl_int_45_27 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c28
+ bl_int_46_28 bl_int_45_28 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c29
+ bl_int_46_29 bl_int_45_29 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c30
+ bl_int_46_30 bl_int_45_30 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c31
+ bl_int_46_31 bl_int_45_31 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c32
+ bl_int_46_32 bl_int_45_32 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c33
+ bl_int_46_33 bl_int_45_33 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c34
+ bl_int_46_34 bl_int_45_34 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c35
+ bl_int_46_35 bl_int_45_35 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c36
+ bl_int_46_36 bl_int_45_36 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c37
+ bl_int_46_37 bl_int_45_37 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c38
+ bl_int_46_38 bl_int_45_38 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c39
+ bl_int_46_39 bl_int_45_39 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c40
+ bl_int_46_40 bl_int_45_40 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c41
+ bl_int_46_41 bl_int_45_41 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c42
+ bl_int_46_42 bl_int_45_42 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c43
+ bl_int_46_43 bl_int_45_43 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c44
+ bl_int_46_44 bl_int_45_44 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c45
+ bl_int_46_45 bl_int_45_45 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c46
+ bl_int_46_46 bl_int_45_46 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c47
+ bl_int_46_47 bl_int_45_47 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c48
+ bl_int_46_48 bl_int_45_48 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c49
+ bl_int_46_49 bl_int_45_49 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c50
+ bl_int_46_50 bl_int_45_50 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c51
+ bl_int_46_51 bl_int_45_51 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c52
+ bl_int_46_52 bl_int_45_52 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c53
+ bl_int_46_53 bl_int_45_53 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c54
+ bl_int_46_54 bl_int_45_54 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c55
+ bl_int_46_55 bl_int_45_55 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c56
+ bl_int_46_56 bl_int_45_56 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c57
+ bl_int_46_57 bl_int_45_57 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c58
+ bl_int_46_58 bl_int_45_58 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c59
+ bl_int_46_59 bl_int_45_59 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c60
+ bl_int_46_60 bl_int_45_60 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c61
+ bl_int_46_61 bl_int_45_61 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c62
+ bl_int_46_62 bl_int_45_62 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c63
+ bl_int_46_63 bl_int_45_63 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c64
+ bl_int_46_64 bl_int_45_64 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c65
+ bl_int_46_65 bl_int_45_65 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c66
+ bl_int_46_66 bl_int_45_66 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c67
+ bl_int_46_67 bl_int_45_67 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c68
+ bl_int_46_68 bl_int_45_68 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c69
+ bl_int_46_69 bl_int_45_69 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c70
+ bl_int_46_70 bl_int_45_70 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c71
+ bl_int_46_71 bl_int_45_71 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c72
+ bl_int_46_72 bl_int_45_72 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c73
+ bl_int_46_73 bl_int_45_73 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c74
+ bl_int_46_74 bl_int_45_74 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c75
+ bl_int_46_75 bl_int_45_75 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c76
+ bl_int_46_76 bl_int_45_76 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c77
+ bl_int_46_77 bl_int_45_77 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c78
+ bl_int_46_78 bl_int_45_78 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c79
+ bl_int_46_79 bl_int_45_79 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c80
+ bl_int_46_80 bl_int_45_80 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c81
+ bl_int_46_81 bl_int_45_81 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c82
+ bl_int_46_82 bl_int_45_82 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c83
+ bl_int_46_83 bl_int_45_83 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c84
+ bl_int_46_84 bl_int_45_84 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c85
+ bl_int_46_85 bl_int_45_85 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c86
+ bl_int_46_86 bl_int_45_86 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c87
+ bl_int_46_87 bl_int_45_87 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c88
+ bl_int_46_88 bl_int_45_88 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c89
+ bl_int_46_89 bl_int_45_89 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c90
+ bl_int_46_90 bl_int_45_90 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c91
+ bl_int_46_91 bl_int_45_91 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c92
+ bl_int_46_92 bl_int_45_92 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c93
+ bl_int_46_93 bl_int_45_93 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c94
+ bl_int_46_94 bl_int_45_94 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c95
+ bl_int_46_95 bl_int_45_95 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c96
+ bl_int_46_96 bl_int_45_96 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c97
+ bl_int_46_97 bl_int_45_97 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c98
+ bl_int_46_98 bl_int_45_98 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c99
+ bl_int_46_99 bl_int_45_99 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c100
+ bl_int_46_100 bl_int_45_100 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c101
+ bl_int_46_101 bl_int_45_101 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c102
+ bl_int_46_102 bl_int_45_102 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c103
+ bl_int_46_103 bl_int_45_103 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c104
+ bl_int_46_104 bl_int_45_104 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c105
+ bl_int_46_105 bl_int_45_105 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c106
+ bl_int_46_106 bl_int_45_106 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c107
+ bl_int_46_107 bl_int_45_107 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c108
+ bl_int_46_108 bl_int_45_108 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c109
+ bl_int_46_109 bl_int_45_109 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c110
+ bl_int_46_110 bl_int_45_110 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c111
+ bl_int_46_111 bl_int_45_111 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c112
+ bl_int_46_112 bl_int_45_112 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c113
+ bl_int_46_113 bl_int_45_113 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c114
+ bl_int_46_114 bl_int_45_114 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c115
+ bl_int_46_115 bl_int_45_115 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c116
+ bl_int_46_116 bl_int_45_116 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c117
+ bl_int_46_117 bl_int_45_117 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c118
+ bl_int_46_118 bl_int_45_118 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c119
+ bl_int_46_119 bl_int_45_119 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c120
+ bl_int_46_120 bl_int_45_120 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c121
+ bl_int_46_121 bl_int_45_121 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c122
+ bl_int_46_122 bl_int_45_122 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c123
+ bl_int_46_123 bl_int_45_123 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c124
+ bl_int_46_124 bl_int_45_124 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c125
+ bl_int_46_125 bl_int_45_125 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c126
+ bl_int_46_126 bl_int_45_126 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c127
+ bl_int_46_127 bl_int_45_127 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c128
+ bl_int_46_128 bl_int_45_128 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c129
+ bl_int_46_129 bl_int_45_129 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c130
+ bl_int_46_130 bl_int_45_130 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c131
+ bl_int_46_131 bl_int_45_131 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c132
+ bl_int_46_132 bl_int_45_132 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c133
+ bl_int_46_133 bl_int_45_133 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c134
+ bl_int_46_134 bl_int_45_134 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c135
+ bl_int_46_135 bl_int_45_135 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c136
+ bl_int_46_136 bl_int_45_136 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c137
+ bl_int_46_137 bl_int_45_137 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c138
+ bl_int_46_138 bl_int_45_138 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c139
+ bl_int_46_139 bl_int_45_139 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c140
+ bl_int_46_140 bl_int_45_140 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c141
+ bl_int_46_141 bl_int_45_141 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c142
+ bl_int_46_142 bl_int_45_142 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c143
+ bl_int_46_143 bl_int_45_143 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c144
+ bl_int_46_144 bl_int_45_144 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c145
+ bl_int_46_145 bl_int_45_145 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c146
+ bl_int_46_146 bl_int_45_146 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c147
+ bl_int_46_147 bl_int_45_147 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c148
+ bl_int_46_148 bl_int_45_148 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c149
+ bl_int_46_149 bl_int_45_149 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c150
+ bl_int_46_150 bl_int_45_150 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c151
+ bl_int_46_151 bl_int_45_151 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c152
+ bl_int_46_152 bl_int_45_152 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c153
+ bl_int_46_153 bl_int_45_153 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c154
+ bl_int_46_154 bl_int_45_154 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c155
+ bl_int_46_155 bl_int_45_155 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c156
+ bl_int_46_156 bl_int_45_156 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c157
+ bl_int_46_157 bl_int_45_157 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c158
+ bl_int_46_158 bl_int_45_158 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c159
+ bl_int_46_159 bl_int_45_159 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c160
+ bl_int_46_160 bl_int_45_160 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c161
+ bl_int_46_161 bl_int_45_161 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c162
+ bl_int_46_162 bl_int_45_162 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c163
+ bl_int_46_163 bl_int_45_163 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c164
+ bl_int_46_164 bl_int_45_164 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c165
+ bl_int_46_165 bl_int_45_165 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c166
+ bl_int_46_166 bl_int_45_166 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c167
+ bl_int_46_167 bl_int_45_167 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c168
+ bl_int_46_168 bl_int_45_168 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c169
+ bl_int_46_169 bl_int_45_169 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c170
+ bl_int_46_170 bl_int_45_170 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c171
+ bl_int_46_171 bl_int_45_171 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c172
+ bl_int_46_172 bl_int_45_172 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c173
+ bl_int_46_173 bl_int_45_173 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c174
+ bl_int_46_174 bl_int_45_174 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c175
+ bl_int_46_175 bl_int_45_175 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c176
+ bl_int_46_176 bl_int_45_176 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c177
+ bl_int_46_177 bl_int_45_177 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c178
+ bl_int_46_178 bl_int_45_178 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c179
+ bl_int_46_179 bl_int_45_179 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c180
+ bl_int_46_180 bl_int_45_180 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c181
+ bl_int_46_181 bl_int_45_181 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c182
+ bl_int_46_182 bl_int_45_182 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r46_c183
+ bl_int_46_183 bl_int_45_183 wl_0_46 gnd
+ sram_rom_base_one_cell
Xbit_r47_c0
+ bl_int_47_0 bl_int_46_0 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c1
+ bl_int_47_1 bl_int_46_1 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c2
+ bl_int_47_2 bl_int_46_2 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c3
+ bl_int_47_3 bl_int_46_3 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c4
+ bl_int_47_4 bl_int_46_4 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c5
+ bl_int_47_5 bl_int_46_5 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c6
+ bl_int_47_6 bl_int_46_6 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c7
+ bl_int_47_7 bl_int_46_7 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c8
+ bl_int_47_8 bl_int_46_8 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c9
+ bl_int_47_9 bl_int_46_9 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c10
+ bl_int_47_10 bl_int_46_10 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c11
+ bl_int_47_11 bl_int_46_11 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c12
+ bl_int_47_12 bl_int_46_12 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c13
+ bl_int_47_13 bl_int_46_13 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c14
+ bl_int_47_14 bl_int_46_14 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c15
+ bl_int_47_15 bl_int_46_15 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c16
+ bl_int_47_16 bl_int_46_16 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c17
+ bl_int_47_17 bl_int_46_17 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c18
+ bl_int_47_18 bl_int_46_18 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c19
+ bl_int_47_19 bl_int_46_19 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c20
+ bl_int_47_20 bl_int_46_20 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c21
+ bl_int_47_21 bl_int_46_21 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c22
+ bl_int_47_22 bl_int_46_22 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c23
+ bl_int_47_23 bl_int_46_23 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c24
+ bl_int_47_24 bl_int_46_24 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c25
+ bl_int_47_25 bl_int_46_25 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c26
+ bl_int_47_26 bl_int_46_26 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c27
+ bl_int_47_27 bl_int_46_27 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c28
+ bl_int_47_28 bl_int_46_28 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c29
+ bl_int_47_29 bl_int_46_29 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c30
+ bl_int_47_30 bl_int_46_30 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c31
+ bl_int_47_31 bl_int_46_31 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c32
+ bl_int_47_32 bl_int_46_32 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c33
+ bl_int_47_33 bl_int_46_33 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c34
+ bl_int_47_34 bl_int_46_34 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c35
+ bl_int_47_35 bl_int_46_35 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c36
+ bl_int_47_36 bl_int_46_36 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c37
+ bl_int_47_37 bl_int_46_37 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c38
+ bl_int_47_38 bl_int_46_38 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c39
+ bl_int_47_39 bl_int_46_39 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c40
+ bl_int_47_40 bl_int_46_40 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c41
+ bl_int_47_41 bl_int_46_41 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c42
+ bl_int_47_42 bl_int_46_42 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c43
+ bl_int_47_43 bl_int_46_43 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c44
+ bl_int_47_44 bl_int_46_44 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c45
+ bl_int_47_45 bl_int_46_45 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c46
+ bl_int_47_46 bl_int_46_46 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c47
+ bl_int_47_47 bl_int_46_47 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c48
+ bl_int_47_48 bl_int_46_48 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c49
+ bl_int_47_49 bl_int_46_49 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c50
+ bl_int_47_50 bl_int_46_50 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c51
+ bl_int_47_51 bl_int_46_51 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c52
+ bl_int_47_52 bl_int_46_52 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c53
+ bl_int_47_53 bl_int_46_53 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c54
+ bl_int_47_54 bl_int_46_54 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c55
+ bl_int_47_55 bl_int_46_55 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c56
+ bl_int_47_56 bl_int_46_56 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c57
+ bl_int_47_57 bl_int_46_57 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c58
+ bl_int_47_58 bl_int_46_58 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c59
+ bl_int_47_59 bl_int_46_59 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c60
+ bl_int_47_60 bl_int_46_60 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c61
+ bl_int_47_61 bl_int_46_61 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c62
+ bl_int_47_62 bl_int_46_62 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c63
+ bl_int_47_63 bl_int_46_63 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c64
+ bl_int_47_64 bl_int_46_64 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c65
+ bl_int_47_65 bl_int_46_65 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c66
+ bl_int_47_66 bl_int_46_66 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c67
+ bl_int_47_67 bl_int_46_67 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c68
+ bl_int_47_68 bl_int_46_68 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c69
+ bl_int_47_69 bl_int_46_69 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c70
+ bl_int_47_70 bl_int_46_70 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c71
+ bl_int_47_71 bl_int_46_71 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c72
+ bl_int_47_72 bl_int_46_72 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c73
+ bl_int_47_73 bl_int_46_73 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c74
+ bl_int_47_74 bl_int_46_74 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c75
+ bl_int_47_75 bl_int_46_75 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c76
+ bl_int_47_76 bl_int_46_76 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c77
+ bl_int_47_77 bl_int_46_77 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c78
+ bl_int_47_78 bl_int_46_78 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c79
+ bl_int_47_79 bl_int_46_79 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c80
+ bl_int_47_80 bl_int_46_80 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c81
+ bl_int_47_81 bl_int_46_81 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c82
+ bl_int_47_82 bl_int_46_82 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c83
+ bl_int_47_83 bl_int_46_83 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c84
+ bl_int_47_84 bl_int_46_84 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c85
+ bl_int_47_85 bl_int_46_85 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c86
+ bl_int_47_86 bl_int_46_86 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c87
+ bl_int_47_87 bl_int_46_87 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c88
+ bl_int_47_88 bl_int_46_88 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c89
+ bl_int_47_89 bl_int_46_89 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c90
+ bl_int_47_90 bl_int_46_90 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c91
+ bl_int_47_91 bl_int_46_91 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c92
+ bl_int_47_92 bl_int_46_92 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c93
+ bl_int_47_93 bl_int_46_93 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c94
+ bl_int_47_94 bl_int_46_94 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c95
+ bl_int_47_95 bl_int_46_95 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c96
+ bl_int_47_96 bl_int_46_96 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c97
+ bl_int_47_97 bl_int_46_97 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c98
+ bl_int_47_98 bl_int_46_98 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c99
+ bl_int_47_99 bl_int_46_99 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c100
+ bl_int_47_100 bl_int_46_100 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c101
+ bl_int_47_101 bl_int_46_101 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c102
+ bl_int_47_102 bl_int_46_102 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c103
+ bl_int_47_103 bl_int_46_103 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c104
+ bl_int_47_104 bl_int_46_104 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c105
+ bl_int_47_105 bl_int_46_105 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c106
+ bl_int_47_106 bl_int_46_106 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c107
+ bl_int_47_107 bl_int_46_107 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c108
+ bl_int_47_108 bl_int_46_108 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c109
+ bl_int_47_109 bl_int_46_109 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c110
+ bl_int_47_110 bl_int_46_110 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c111
+ bl_int_47_111 bl_int_46_111 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c112
+ bl_int_47_112 bl_int_46_112 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c113
+ bl_int_47_113 bl_int_46_113 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c114
+ bl_int_47_114 bl_int_46_114 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c115
+ bl_int_47_115 bl_int_46_115 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c116
+ bl_int_47_116 bl_int_46_116 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c117
+ bl_int_47_117 bl_int_46_117 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c118
+ bl_int_47_118 bl_int_46_118 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c119
+ bl_int_47_119 bl_int_46_119 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c120
+ bl_int_47_120 bl_int_46_120 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c121
+ bl_int_47_121 bl_int_46_121 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c122
+ bl_int_47_122 bl_int_46_122 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c123
+ bl_int_47_123 bl_int_46_123 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c124
+ bl_int_47_124 bl_int_46_124 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c125
+ bl_int_47_125 bl_int_46_125 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c126
+ bl_int_47_126 bl_int_46_126 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c127
+ bl_int_47_127 bl_int_46_127 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c128
+ bl_int_47_128 bl_int_46_128 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c129
+ bl_int_47_129 bl_int_46_129 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c130
+ bl_int_47_130 bl_int_46_130 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c131
+ bl_int_47_131 bl_int_46_131 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c132
+ bl_int_47_132 bl_int_46_132 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c133
+ bl_int_47_133 bl_int_46_133 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c134
+ bl_int_47_134 bl_int_46_134 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c135
+ bl_int_47_135 bl_int_46_135 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c136
+ bl_int_47_136 bl_int_46_136 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c137
+ bl_int_47_137 bl_int_46_137 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c138
+ bl_int_47_138 bl_int_46_138 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c139
+ bl_int_47_139 bl_int_46_139 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c140
+ bl_int_47_140 bl_int_46_140 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c141
+ bl_int_47_141 bl_int_46_141 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c142
+ bl_int_47_142 bl_int_46_142 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c143
+ bl_int_47_143 bl_int_46_143 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c144
+ bl_int_47_144 bl_int_46_144 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c145
+ bl_int_47_145 bl_int_46_145 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c146
+ bl_int_47_146 bl_int_46_146 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c147
+ bl_int_47_147 bl_int_46_147 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c148
+ bl_int_47_148 bl_int_46_148 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c149
+ bl_int_47_149 bl_int_46_149 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c150
+ bl_int_47_150 bl_int_46_150 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c151
+ bl_int_47_151 bl_int_46_151 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c152
+ bl_int_47_152 bl_int_46_152 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c153
+ bl_int_47_153 bl_int_46_153 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c154
+ bl_int_47_154 bl_int_46_154 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c155
+ bl_int_47_155 bl_int_46_155 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c156
+ bl_int_47_156 bl_int_46_156 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c157
+ bl_int_47_157 bl_int_46_157 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c158
+ bl_int_47_158 bl_int_46_158 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c159
+ bl_int_47_159 bl_int_46_159 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c160
+ bl_int_47_160 bl_int_46_160 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c161
+ bl_int_47_161 bl_int_46_161 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c162
+ bl_int_47_162 bl_int_46_162 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c163
+ bl_int_47_163 bl_int_46_163 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c164
+ bl_int_47_164 bl_int_46_164 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c165
+ bl_int_47_165 bl_int_46_165 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c166
+ bl_int_47_166 bl_int_46_166 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c167
+ bl_int_47_167 bl_int_46_167 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c168
+ bl_int_47_168 bl_int_46_168 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c169
+ bl_int_47_169 bl_int_46_169 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c170
+ bl_int_47_170 bl_int_46_170 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c171
+ bl_int_47_171 bl_int_46_171 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c172
+ bl_int_47_172 bl_int_46_172 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c173
+ bl_int_47_173 bl_int_46_173 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c174
+ bl_int_47_174 bl_int_46_174 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c175
+ bl_int_47_175 bl_int_46_175 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c176
+ bl_int_47_176 bl_int_46_176 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c177
+ bl_int_47_177 bl_int_46_177 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c178
+ bl_int_47_178 bl_int_46_178 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c179
+ bl_int_47_179 bl_int_46_179 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c180
+ bl_int_47_180 bl_int_46_180 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c181
+ bl_int_47_181 bl_int_46_181 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c182
+ bl_int_47_182 bl_int_46_182 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r47_c183
+ bl_int_47_183 bl_int_46_183 wl_0_47 gnd
+ sram_rom_base_one_cell
Xbit_r48_c0
+ bl_int_48_0 bl_int_47_0 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c1
+ bl_int_48_1 bl_int_47_1 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c2
+ bl_int_48_2 bl_int_47_2 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c3
+ bl_int_48_3 bl_int_47_3 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c4
+ bl_int_48_4 bl_int_47_4 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c5
+ bl_int_48_5 bl_int_47_5 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c6
+ bl_int_48_6 bl_int_47_6 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c7
+ bl_int_48_7 bl_int_47_7 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c8
+ bl_int_48_8 bl_int_47_8 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c9
+ bl_int_48_9 bl_int_47_9 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c10
+ bl_int_48_10 bl_int_47_10 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c11
+ bl_int_48_11 bl_int_47_11 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c12
+ bl_int_48_12 bl_int_47_12 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c13
+ bl_int_48_13 bl_int_47_13 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c14
+ bl_int_48_14 bl_int_47_14 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c15
+ bl_int_48_15 bl_int_47_15 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c16
+ bl_int_48_16 bl_int_47_16 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c17
+ bl_int_48_17 bl_int_47_17 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c18
+ bl_int_48_18 bl_int_47_18 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c19
+ bl_int_48_19 bl_int_47_19 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c20
+ bl_int_48_20 bl_int_47_20 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c21
+ bl_int_48_21 bl_int_47_21 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c22
+ bl_int_48_22 bl_int_47_22 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c23
+ bl_int_48_23 bl_int_47_23 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c24
+ bl_int_48_24 bl_int_47_24 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c25
+ bl_int_48_25 bl_int_47_25 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c26
+ bl_int_48_26 bl_int_47_26 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c27
+ bl_int_48_27 bl_int_47_27 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c28
+ bl_int_48_28 bl_int_47_28 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c29
+ bl_int_48_29 bl_int_47_29 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c30
+ bl_int_48_30 bl_int_47_30 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c31
+ bl_int_48_31 bl_int_47_31 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c32
+ bl_int_48_32 bl_int_47_32 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c33
+ bl_int_48_33 bl_int_47_33 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c34
+ bl_int_48_34 bl_int_47_34 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c35
+ bl_int_48_35 bl_int_47_35 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c36
+ bl_int_48_36 bl_int_47_36 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c37
+ bl_int_48_37 bl_int_47_37 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c38
+ bl_int_48_38 bl_int_47_38 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c39
+ bl_int_48_39 bl_int_47_39 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c40
+ bl_int_48_40 bl_int_47_40 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c41
+ bl_int_48_41 bl_int_47_41 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c42
+ bl_int_48_42 bl_int_47_42 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c43
+ bl_int_48_43 bl_int_47_43 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c44
+ bl_int_48_44 bl_int_47_44 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c45
+ bl_int_48_45 bl_int_47_45 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c46
+ bl_int_48_46 bl_int_47_46 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c47
+ bl_int_48_47 bl_int_47_47 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c48
+ bl_int_48_48 bl_int_47_48 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c49
+ bl_int_48_49 bl_int_47_49 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c50
+ bl_int_48_50 bl_int_47_50 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c51
+ bl_int_48_51 bl_int_47_51 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c52
+ bl_int_48_52 bl_int_47_52 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c53
+ bl_int_48_53 bl_int_47_53 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c54
+ bl_int_48_54 bl_int_47_54 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c55
+ bl_int_48_55 bl_int_47_55 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c56
+ bl_int_48_56 bl_int_47_56 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c57
+ bl_int_48_57 bl_int_47_57 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c58
+ bl_int_48_58 bl_int_47_58 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c59
+ bl_int_48_59 bl_int_47_59 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c60
+ bl_int_48_60 bl_int_47_60 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c61
+ bl_int_48_61 bl_int_47_61 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c62
+ bl_int_48_62 bl_int_47_62 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c63
+ bl_int_48_63 bl_int_47_63 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c64
+ bl_int_48_64 bl_int_47_64 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c65
+ bl_int_48_65 bl_int_47_65 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c66
+ bl_int_48_66 bl_int_47_66 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c67
+ bl_int_48_67 bl_int_47_67 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c68
+ bl_int_48_68 bl_int_47_68 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c69
+ bl_int_48_69 bl_int_47_69 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c70
+ bl_int_48_70 bl_int_47_70 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c71
+ bl_int_48_71 bl_int_47_71 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c72
+ bl_int_48_72 bl_int_47_72 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c73
+ bl_int_48_73 bl_int_47_73 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c74
+ bl_int_48_74 bl_int_47_74 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c75
+ bl_int_48_75 bl_int_47_75 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c76
+ bl_int_48_76 bl_int_47_76 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c77
+ bl_int_48_77 bl_int_47_77 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c78
+ bl_int_48_78 bl_int_47_78 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c79
+ bl_int_48_79 bl_int_47_79 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c80
+ bl_int_48_80 bl_int_47_80 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c81
+ bl_int_48_81 bl_int_47_81 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c82
+ bl_int_48_82 bl_int_47_82 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c83
+ bl_int_48_83 bl_int_47_83 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c84
+ bl_int_48_84 bl_int_47_84 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c85
+ bl_int_48_85 bl_int_47_85 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c86
+ bl_int_48_86 bl_int_47_86 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c87
+ bl_int_48_87 bl_int_47_87 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c88
+ bl_int_48_88 bl_int_47_88 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c89
+ bl_int_48_89 bl_int_47_89 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c90
+ bl_int_48_90 bl_int_47_90 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c91
+ bl_int_48_91 bl_int_47_91 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c92
+ bl_int_48_92 bl_int_47_92 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c93
+ bl_int_48_93 bl_int_47_93 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c94
+ bl_int_48_94 bl_int_47_94 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c95
+ bl_int_48_95 bl_int_47_95 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c96
+ bl_int_48_96 bl_int_47_96 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c97
+ bl_int_48_97 bl_int_47_97 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c98
+ bl_int_48_98 bl_int_47_98 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c99
+ bl_int_48_99 bl_int_47_99 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c100
+ bl_int_48_100 bl_int_47_100 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c101
+ bl_int_48_101 bl_int_47_101 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c102
+ bl_int_48_102 bl_int_47_102 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c103
+ bl_int_48_103 bl_int_47_103 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c104
+ bl_int_48_104 bl_int_47_104 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c105
+ bl_int_48_105 bl_int_47_105 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c106
+ bl_int_48_106 bl_int_47_106 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c107
+ bl_int_48_107 bl_int_47_107 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c108
+ bl_int_48_108 bl_int_47_108 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c109
+ bl_int_48_109 bl_int_47_109 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c110
+ bl_int_48_110 bl_int_47_110 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c111
+ bl_int_48_111 bl_int_47_111 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c112
+ bl_int_48_112 bl_int_47_112 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c113
+ bl_int_48_113 bl_int_47_113 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c114
+ bl_int_48_114 bl_int_47_114 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c115
+ bl_int_48_115 bl_int_47_115 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c116
+ bl_int_48_116 bl_int_47_116 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c117
+ bl_int_48_117 bl_int_47_117 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c118
+ bl_int_48_118 bl_int_47_118 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c119
+ bl_int_48_119 bl_int_47_119 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c120
+ bl_int_48_120 bl_int_47_120 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c121
+ bl_int_48_121 bl_int_47_121 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c122
+ bl_int_48_122 bl_int_47_122 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c123
+ bl_int_48_123 bl_int_47_123 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c124
+ bl_int_48_124 bl_int_47_124 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c125
+ bl_int_48_125 bl_int_47_125 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c126
+ bl_int_48_126 bl_int_47_126 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c127
+ bl_int_48_127 bl_int_47_127 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c128
+ bl_int_48_128 bl_int_47_128 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c129
+ bl_int_48_129 bl_int_47_129 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c130
+ bl_int_48_130 bl_int_47_130 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c131
+ bl_int_48_131 bl_int_47_131 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c132
+ bl_int_48_132 bl_int_47_132 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c133
+ bl_int_48_133 bl_int_47_133 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c134
+ bl_int_48_134 bl_int_47_134 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c135
+ bl_int_48_135 bl_int_47_135 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c136
+ bl_int_48_136 bl_int_47_136 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c137
+ bl_int_48_137 bl_int_47_137 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c138
+ bl_int_48_138 bl_int_47_138 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c139
+ bl_int_48_139 bl_int_47_139 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c140
+ bl_int_48_140 bl_int_47_140 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c141
+ bl_int_48_141 bl_int_47_141 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c142
+ bl_int_48_142 bl_int_47_142 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c143
+ bl_int_48_143 bl_int_47_143 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c144
+ bl_int_48_144 bl_int_47_144 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c145
+ bl_int_48_145 bl_int_47_145 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c146
+ bl_int_48_146 bl_int_47_146 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c147
+ bl_int_48_147 bl_int_47_147 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c148
+ bl_int_48_148 bl_int_47_148 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c149
+ bl_int_48_149 bl_int_47_149 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c150
+ bl_int_48_150 bl_int_47_150 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c151
+ bl_int_48_151 bl_int_47_151 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c152
+ bl_int_48_152 bl_int_47_152 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c153
+ bl_int_48_153 bl_int_47_153 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c154
+ bl_int_48_154 bl_int_47_154 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c155
+ bl_int_48_155 bl_int_47_155 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c156
+ bl_int_48_156 bl_int_47_156 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c157
+ bl_int_48_157 bl_int_47_157 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c158
+ bl_int_48_158 bl_int_47_158 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c159
+ bl_int_48_159 bl_int_47_159 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c160
+ bl_int_48_160 bl_int_47_160 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c161
+ bl_int_48_161 bl_int_47_161 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c162
+ bl_int_48_162 bl_int_47_162 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c163
+ bl_int_48_163 bl_int_47_163 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c164
+ bl_int_48_164 bl_int_47_164 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c165
+ bl_int_48_165 bl_int_47_165 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c166
+ bl_int_48_166 bl_int_47_166 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c167
+ bl_int_48_167 bl_int_47_167 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c168
+ bl_int_48_168 bl_int_47_168 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c169
+ bl_int_48_169 bl_int_47_169 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c170
+ bl_int_48_170 bl_int_47_170 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c171
+ bl_int_48_171 bl_int_47_171 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c172
+ bl_int_48_172 bl_int_47_172 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c173
+ bl_int_48_173 bl_int_47_173 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c174
+ bl_int_48_174 bl_int_47_174 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c175
+ bl_int_48_175 bl_int_47_175 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c176
+ bl_int_48_176 bl_int_47_176 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c177
+ bl_int_48_177 bl_int_47_177 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c178
+ bl_int_48_178 bl_int_47_178 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c179
+ bl_int_48_179 bl_int_47_179 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c180
+ bl_int_48_180 bl_int_47_180 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c181
+ bl_int_48_181 bl_int_47_181 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c182
+ bl_int_48_182 bl_int_47_182 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r48_c183
+ bl_int_48_183 bl_int_47_183 wl_0_48 gnd
+ sram_rom_base_one_cell
Xbit_r49_c0
+ bl_int_49_0 bl_int_48_0 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c1
+ bl_int_49_1 bl_int_48_1 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c2
+ bl_int_49_2 bl_int_48_2 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c3
+ bl_int_49_3 bl_int_48_3 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c4
+ bl_int_49_4 bl_int_48_4 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c5
+ bl_int_49_5 bl_int_48_5 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c6
+ bl_int_49_6 bl_int_48_6 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c7
+ bl_int_49_7 bl_int_48_7 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c8
+ bl_int_49_8 bl_int_48_8 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c9
+ bl_int_49_9 bl_int_48_9 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c10
+ bl_int_49_10 bl_int_48_10 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c11
+ bl_int_49_11 bl_int_48_11 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c12
+ bl_int_49_12 bl_int_48_12 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c13
+ bl_int_49_13 bl_int_48_13 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c14
+ bl_int_49_14 bl_int_48_14 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c15
+ bl_int_49_15 bl_int_48_15 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c16
+ bl_int_49_16 bl_int_48_16 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c17
+ bl_int_49_17 bl_int_48_17 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c18
+ bl_int_49_18 bl_int_48_18 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c19
+ bl_int_49_19 bl_int_48_19 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c20
+ bl_int_49_20 bl_int_48_20 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c21
+ bl_int_49_21 bl_int_48_21 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c22
+ bl_int_49_22 bl_int_48_22 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c23
+ bl_int_49_23 bl_int_48_23 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c24
+ bl_int_49_24 bl_int_48_24 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c25
+ bl_int_49_25 bl_int_48_25 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c26
+ bl_int_49_26 bl_int_48_26 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c27
+ bl_int_49_27 bl_int_48_27 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c28
+ bl_int_49_28 bl_int_48_28 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c29
+ bl_int_49_29 bl_int_48_29 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c30
+ bl_int_49_30 bl_int_48_30 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c31
+ bl_int_49_31 bl_int_48_31 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c32
+ bl_int_49_32 bl_int_48_32 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c33
+ bl_int_49_33 bl_int_48_33 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c34
+ bl_int_49_34 bl_int_48_34 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c35
+ bl_int_49_35 bl_int_48_35 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c36
+ bl_int_49_36 bl_int_48_36 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c37
+ bl_int_49_37 bl_int_48_37 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c38
+ bl_int_49_38 bl_int_48_38 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c39
+ bl_int_49_39 bl_int_48_39 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c40
+ bl_int_49_40 bl_int_48_40 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c41
+ bl_int_49_41 bl_int_48_41 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c42
+ bl_int_49_42 bl_int_48_42 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c43
+ bl_int_49_43 bl_int_48_43 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c44
+ bl_int_49_44 bl_int_48_44 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c45
+ bl_int_49_45 bl_int_48_45 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c46
+ bl_int_49_46 bl_int_48_46 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c47
+ bl_int_49_47 bl_int_48_47 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c48
+ bl_int_49_48 bl_int_48_48 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c49
+ bl_int_49_49 bl_int_48_49 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c50
+ bl_int_49_50 bl_int_48_50 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c51
+ bl_int_49_51 bl_int_48_51 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c52
+ bl_int_49_52 bl_int_48_52 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c53
+ bl_int_49_53 bl_int_48_53 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c54
+ bl_int_49_54 bl_int_48_54 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c55
+ bl_int_49_55 bl_int_48_55 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c56
+ bl_int_49_56 bl_int_48_56 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c57
+ bl_int_49_57 bl_int_48_57 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c58
+ bl_int_49_58 bl_int_48_58 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c59
+ bl_int_49_59 bl_int_48_59 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c60
+ bl_int_49_60 bl_int_48_60 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c61
+ bl_int_49_61 bl_int_48_61 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c62
+ bl_int_49_62 bl_int_48_62 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c63
+ bl_int_49_63 bl_int_48_63 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c64
+ bl_int_49_64 bl_int_48_64 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c65
+ bl_int_49_65 bl_int_48_65 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c66
+ bl_int_49_66 bl_int_48_66 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c67
+ bl_int_49_67 bl_int_48_67 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c68
+ bl_int_49_68 bl_int_48_68 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c69
+ bl_int_49_69 bl_int_48_69 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c70
+ bl_int_49_70 bl_int_48_70 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c71
+ bl_int_49_71 bl_int_48_71 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c72
+ bl_int_49_72 bl_int_48_72 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c73
+ bl_int_49_73 bl_int_48_73 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c74
+ bl_int_49_74 bl_int_48_74 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c75
+ bl_int_49_75 bl_int_48_75 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c76
+ bl_int_49_76 bl_int_48_76 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c77
+ bl_int_49_77 bl_int_48_77 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c78
+ bl_int_49_78 bl_int_48_78 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c79
+ bl_int_49_79 bl_int_48_79 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c80
+ bl_int_49_80 bl_int_48_80 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c81
+ bl_int_49_81 bl_int_48_81 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c82
+ bl_int_49_82 bl_int_48_82 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c83
+ bl_int_49_83 bl_int_48_83 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c84
+ bl_int_49_84 bl_int_48_84 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c85
+ bl_int_49_85 bl_int_48_85 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c86
+ bl_int_49_86 bl_int_48_86 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c87
+ bl_int_49_87 bl_int_48_87 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c88
+ bl_int_49_88 bl_int_48_88 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c89
+ bl_int_49_89 bl_int_48_89 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c90
+ bl_int_49_90 bl_int_48_90 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c91
+ bl_int_49_91 bl_int_48_91 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c92
+ bl_int_49_92 bl_int_48_92 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c93
+ bl_int_49_93 bl_int_48_93 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c94
+ bl_int_49_94 bl_int_48_94 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c95
+ bl_int_49_95 bl_int_48_95 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c96
+ bl_int_49_96 bl_int_48_96 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c97
+ bl_int_49_97 bl_int_48_97 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c98
+ bl_int_49_98 bl_int_48_98 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c99
+ bl_int_49_99 bl_int_48_99 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c100
+ bl_int_49_100 bl_int_48_100 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c101
+ bl_int_49_101 bl_int_48_101 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c102
+ bl_int_49_102 bl_int_48_102 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c103
+ bl_int_49_103 bl_int_48_103 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c104
+ bl_int_49_104 bl_int_48_104 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c105
+ bl_int_49_105 bl_int_48_105 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c106
+ bl_int_49_106 bl_int_48_106 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c107
+ bl_int_49_107 bl_int_48_107 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c108
+ bl_int_49_108 bl_int_48_108 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c109
+ bl_int_49_109 bl_int_48_109 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c110
+ bl_int_49_110 bl_int_48_110 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c111
+ bl_int_49_111 bl_int_48_111 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c112
+ bl_int_49_112 bl_int_48_112 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c113
+ bl_int_49_113 bl_int_48_113 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c114
+ bl_int_49_114 bl_int_48_114 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c115
+ bl_int_49_115 bl_int_48_115 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c116
+ bl_int_49_116 bl_int_48_116 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c117
+ bl_int_49_117 bl_int_48_117 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c118
+ bl_int_49_118 bl_int_48_118 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c119
+ bl_int_49_119 bl_int_48_119 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c120
+ bl_int_49_120 bl_int_48_120 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c121
+ bl_int_49_121 bl_int_48_121 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c122
+ bl_int_49_122 bl_int_48_122 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c123
+ bl_int_49_123 bl_int_48_123 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c124
+ bl_int_49_124 bl_int_48_124 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c125
+ bl_int_49_125 bl_int_48_125 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c126
+ bl_int_49_126 bl_int_48_126 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c127
+ bl_int_49_127 bl_int_48_127 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c128
+ bl_int_49_128 bl_int_48_128 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c129
+ bl_int_49_129 bl_int_48_129 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c130
+ bl_int_49_130 bl_int_48_130 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c131
+ bl_int_49_131 bl_int_48_131 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c132
+ bl_int_49_132 bl_int_48_132 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c133
+ bl_int_49_133 bl_int_48_133 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c134
+ bl_int_49_134 bl_int_48_134 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c135
+ bl_int_49_135 bl_int_48_135 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c136
+ bl_int_49_136 bl_int_48_136 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c137
+ bl_int_49_137 bl_int_48_137 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c138
+ bl_int_49_138 bl_int_48_138 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c139
+ bl_int_49_139 bl_int_48_139 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c140
+ bl_int_49_140 bl_int_48_140 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c141
+ bl_int_49_141 bl_int_48_141 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c142
+ bl_int_49_142 bl_int_48_142 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c143
+ bl_int_49_143 bl_int_48_143 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c144
+ bl_int_49_144 bl_int_48_144 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c145
+ bl_int_49_145 bl_int_48_145 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c146
+ bl_int_49_146 bl_int_48_146 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c147
+ bl_int_49_147 bl_int_48_147 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c148
+ bl_int_49_148 bl_int_48_148 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c149
+ bl_int_49_149 bl_int_48_149 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c150
+ bl_int_49_150 bl_int_48_150 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c151
+ bl_int_49_151 bl_int_48_151 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c152
+ bl_int_49_152 bl_int_48_152 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c153
+ bl_int_49_153 bl_int_48_153 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c154
+ bl_int_49_154 bl_int_48_154 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c155
+ bl_int_49_155 bl_int_48_155 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c156
+ bl_int_49_156 bl_int_48_156 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c157
+ bl_int_49_157 bl_int_48_157 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c158
+ bl_int_49_158 bl_int_48_158 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c159
+ bl_int_49_159 bl_int_48_159 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c160
+ bl_int_49_160 bl_int_48_160 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c161
+ bl_int_49_161 bl_int_48_161 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c162
+ bl_int_49_162 bl_int_48_162 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c163
+ bl_int_49_163 bl_int_48_163 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c164
+ bl_int_49_164 bl_int_48_164 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c165
+ bl_int_49_165 bl_int_48_165 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c166
+ bl_int_49_166 bl_int_48_166 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c167
+ bl_int_49_167 bl_int_48_167 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c168
+ bl_int_49_168 bl_int_48_168 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c169
+ bl_int_49_169 bl_int_48_169 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c170
+ bl_int_49_170 bl_int_48_170 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c171
+ bl_int_49_171 bl_int_48_171 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c172
+ bl_int_49_172 bl_int_48_172 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c173
+ bl_int_49_173 bl_int_48_173 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c174
+ bl_int_49_174 bl_int_48_174 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c175
+ bl_int_49_175 bl_int_48_175 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c176
+ bl_int_49_176 bl_int_48_176 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c177
+ bl_int_49_177 bl_int_48_177 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c178
+ bl_int_49_178 bl_int_48_178 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c179
+ bl_int_49_179 bl_int_48_179 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c180
+ bl_int_49_180 bl_int_48_180 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c181
+ bl_int_49_181 bl_int_48_181 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c182
+ bl_int_49_182 bl_int_48_182 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r49_c183
+ bl_int_49_183 bl_int_48_183 wl_0_49 gnd
+ sram_rom_base_one_cell
Xbit_r50_c0
+ bl_int_50_0 bl_int_49_0 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c1
+ bl_int_50_1 bl_int_49_1 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c2
+ bl_int_50_2 bl_int_49_2 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c3
+ bl_int_50_3 bl_int_49_3 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c4
+ bl_int_50_4 bl_int_49_4 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c5
+ bl_int_50_5 bl_int_49_5 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c6
+ bl_int_50_6 bl_int_49_6 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c7
+ bl_int_50_7 bl_int_49_7 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c8
+ bl_int_50_8 bl_int_49_8 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c9
+ bl_int_50_9 bl_int_49_9 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c10
+ bl_int_50_10 bl_int_49_10 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c11
+ bl_int_50_11 bl_int_49_11 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c12
+ bl_int_50_12 bl_int_49_12 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c13
+ bl_int_50_13 bl_int_49_13 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c14
+ bl_int_50_14 bl_int_49_14 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c15
+ bl_int_50_15 bl_int_49_15 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c16
+ bl_int_50_16 bl_int_49_16 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c17
+ bl_int_50_17 bl_int_49_17 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c18
+ bl_int_50_18 bl_int_49_18 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c19
+ bl_int_50_19 bl_int_49_19 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c20
+ bl_int_50_20 bl_int_49_20 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c21
+ bl_int_50_21 bl_int_49_21 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c22
+ bl_int_50_22 bl_int_49_22 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c23
+ bl_int_50_23 bl_int_49_23 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c24
+ bl_int_50_24 bl_int_49_24 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c25
+ bl_int_50_25 bl_int_49_25 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c26
+ bl_int_50_26 bl_int_49_26 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c27
+ bl_int_50_27 bl_int_49_27 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c28
+ bl_int_50_28 bl_int_49_28 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c29
+ bl_int_50_29 bl_int_49_29 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c30
+ bl_int_50_30 bl_int_49_30 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c31
+ bl_int_50_31 bl_int_49_31 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c32
+ bl_int_50_32 bl_int_49_32 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c33
+ bl_int_50_33 bl_int_49_33 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c34
+ bl_int_50_34 bl_int_49_34 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c35
+ bl_int_50_35 bl_int_49_35 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c36
+ bl_int_50_36 bl_int_49_36 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c37
+ bl_int_50_37 bl_int_49_37 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c38
+ bl_int_50_38 bl_int_49_38 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c39
+ bl_int_50_39 bl_int_49_39 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c40
+ bl_int_50_40 bl_int_49_40 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c41
+ bl_int_50_41 bl_int_49_41 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c42
+ bl_int_50_42 bl_int_49_42 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c43
+ bl_int_50_43 bl_int_49_43 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c44
+ bl_int_50_44 bl_int_49_44 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c45
+ bl_int_50_45 bl_int_49_45 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c46
+ bl_int_50_46 bl_int_49_46 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c47
+ bl_int_50_47 bl_int_49_47 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c48
+ bl_int_50_48 bl_int_49_48 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c49
+ bl_int_50_49 bl_int_49_49 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c50
+ bl_int_50_50 bl_int_49_50 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c51
+ bl_int_50_51 bl_int_49_51 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c52
+ bl_int_50_52 bl_int_49_52 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c53
+ bl_int_50_53 bl_int_49_53 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c54
+ bl_int_50_54 bl_int_49_54 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c55
+ bl_int_50_55 bl_int_49_55 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c56
+ bl_int_50_56 bl_int_49_56 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c57
+ bl_int_50_57 bl_int_49_57 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c58
+ bl_int_50_58 bl_int_49_58 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c59
+ bl_int_50_59 bl_int_49_59 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c60
+ bl_int_50_60 bl_int_49_60 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c61
+ bl_int_50_61 bl_int_49_61 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c62
+ bl_int_50_62 bl_int_49_62 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c63
+ bl_int_50_63 bl_int_49_63 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c64
+ bl_int_50_64 bl_int_49_64 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c65
+ bl_int_50_65 bl_int_49_65 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c66
+ bl_int_50_66 bl_int_49_66 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c67
+ bl_int_50_67 bl_int_49_67 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c68
+ bl_int_50_68 bl_int_49_68 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c69
+ bl_int_50_69 bl_int_49_69 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c70
+ bl_int_50_70 bl_int_49_70 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c71
+ bl_int_50_71 bl_int_49_71 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c72
+ bl_int_50_72 bl_int_49_72 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c73
+ bl_int_50_73 bl_int_49_73 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c74
+ bl_int_50_74 bl_int_49_74 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c75
+ bl_int_50_75 bl_int_49_75 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c76
+ bl_int_50_76 bl_int_49_76 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c77
+ bl_int_50_77 bl_int_49_77 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c78
+ bl_int_50_78 bl_int_49_78 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c79
+ bl_int_50_79 bl_int_49_79 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c80
+ bl_int_50_80 bl_int_49_80 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c81
+ bl_int_50_81 bl_int_49_81 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c82
+ bl_int_50_82 bl_int_49_82 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c83
+ bl_int_50_83 bl_int_49_83 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c84
+ bl_int_50_84 bl_int_49_84 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c85
+ bl_int_50_85 bl_int_49_85 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c86
+ bl_int_50_86 bl_int_49_86 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c87
+ bl_int_50_87 bl_int_49_87 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c88
+ bl_int_50_88 bl_int_49_88 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c89
+ bl_int_50_89 bl_int_49_89 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c90
+ bl_int_50_90 bl_int_49_90 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c91
+ bl_int_50_91 bl_int_49_91 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c92
+ bl_int_50_92 bl_int_49_92 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c93
+ bl_int_50_93 bl_int_49_93 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c94
+ bl_int_50_94 bl_int_49_94 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c95
+ bl_int_50_95 bl_int_49_95 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c96
+ bl_int_50_96 bl_int_49_96 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c97
+ bl_int_50_97 bl_int_49_97 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c98
+ bl_int_50_98 bl_int_49_98 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c99
+ bl_int_50_99 bl_int_49_99 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c100
+ bl_int_50_100 bl_int_49_100 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c101
+ bl_int_50_101 bl_int_49_101 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c102
+ bl_int_50_102 bl_int_49_102 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c103
+ bl_int_50_103 bl_int_49_103 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c104
+ bl_int_50_104 bl_int_49_104 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c105
+ bl_int_50_105 bl_int_49_105 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c106
+ bl_int_50_106 bl_int_49_106 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c107
+ bl_int_50_107 bl_int_49_107 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c108
+ bl_int_50_108 bl_int_49_108 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c109
+ bl_int_50_109 bl_int_49_109 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c110
+ bl_int_50_110 bl_int_49_110 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c111
+ bl_int_50_111 bl_int_49_111 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c112
+ bl_int_50_112 bl_int_49_112 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c113
+ bl_int_50_113 bl_int_49_113 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c114
+ bl_int_50_114 bl_int_49_114 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c115
+ bl_int_50_115 bl_int_49_115 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c116
+ bl_int_50_116 bl_int_49_116 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c117
+ bl_int_50_117 bl_int_49_117 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c118
+ bl_int_50_118 bl_int_49_118 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c119
+ bl_int_50_119 bl_int_49_119 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c120
+ bl_int_50_120 bl_int_49_120 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c121
+ bl_int_50_121 bl_int_49_121 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c122
+ bl_int_50_122 bl_int_49_122 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c123
+ bl_int_50_123 bl_int_49_123 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c124
+ bl_int_50_124 bl_int_49_124 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c125
+ bl_int_50_125 bl_int_49_125 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c126
+ bl_int_50_126 bl_int_49_126 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c127
+ bl_int_50_127 bl_int_49_127 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c128
+ bl_int_50_128 bl_int_49_128 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c129
+ bl_int_50_129 bl_int_49_129 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c130
+ bl_int_50_130 bl_int_49_130 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c131
+ bl_int_50_131 bl_int_49_131 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c132
+ bl_int_50_132 bl_int_49_132 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c133
+ bl_int_50_133 bl_int_49_133 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c134
+ bl_int_50_134 bl_int_49_134 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c135
+ bl_int_50_135 bl_int_49_135 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c136
+ bl_int_50_136 bl_int_49_136 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c137
+ bl_int_50_137 bl_int_49_137 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c138
+ bl_int_50_138 bl_int_49_138 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c139
+ bl_int_50_139 bl_int_49_139 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c140
+ bl_int_50_140 bl_int_49_140 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c141
+ bl_int_50_141 bl_int_49_141 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c142
+ bl_int_50_142 bl_int_49_142 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c143
+ bl_int_50_143 bl_int_49_143 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c144
+ bl_int_50_144 bl_int_49_144 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c145
+ bl_int_50_145 bl_int_49_145 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c146
+ bl_int_50_146 bl_int_49_146 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c147
+ bl_int_50_147 bl_int_49_147 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c148
+ bl_int_50_148 bl_int_49_148 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c149
+ bl_int_50_149 bl_int_49_149 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c150
+ bl_int_50_150 bl_int_49_150 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c151
+ bl_int_50_151 bl_int_49_151 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c152
+ bl_int_50_152 bl_int_49_152 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c153
+ bl_int_50_153 bl_int_49_153 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c154
+ bl_int_50_154 bl_int_49_154 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c155
+ bl_int_50_155 bl_int_49_155 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c156
+ bl_int_50_156 bl_int_49_156 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c157
+ bl_int_50_157 bl_int_49_157 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c158
+ bl_int_50_158 bl_int_49_158 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c159
+ bl_int_50_159 bl_int_49_159 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c160
+ bl_int_50_160 bl_int_49_160 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c161
+ bl_int_50_161 bl_int_49_161 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c162
+ bl_int_50_162 bl_int_49_162 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c163
+ bl_int_50_163 bl_int_49_163 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c164
+ bl_int_50_164 bl_int_49_164 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c165
+ bl_int_50_165 bl_int_49_165 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c166
+ bl_int_50_166 bl_int_49_166 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c167
+ bl_int_50_167 bl_int_49_167 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c168
+ bl_int_50_168 bl_int_49_168 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c169
+ bl_int_50_169 bl_int_49_169 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c170
+ bl_int_50_170 bl_int_49_170 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c171
+ bl_int_50_171 bl_int_49_171 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c172
+ bl_int_50_172 bl_int_49_172 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c173
+ bl_int_50_173 bl_int_49_173 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c174
+ bl_int_50_174 bl_int_49_174 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c175
+ bl_int_50_175 bl_int_49_175 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c176
+ bl_int_50_176 bl_int_49_176 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c177
+ bl_int_50_177 bl_int_49_177 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c178
+ bl_int_50_178 bl_int_49_178 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c179
+ bl_int_50_179 bl_int_49_179 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c180
+ bl_int_50_180 bl_int_49_180 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c181
+ bl_int_50_181 bl_int_49_181 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c182
+ bl_int_50_182 bl_int_49_182 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r50_c183
+ bl_int_50_183 bl_int_49_183 wl_0_50 gnd
+ sram_rom_base_one_cell
Xbit_r51_c0
+ bl_int_51_0 bl_int_50_0 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c1
+ bl_int_51_1 bl_int_50_1 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c2
+ bl_int_51_2 bl_int_50_2 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c3
+ bl_int_51_3 bl_int_50_3 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c4
+ bl_int_51_4 bl_int_50_4 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c5
+ bl_int_51_5 bl_int_50_5 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c6
+ bl_int_51_6 bl_int_50_6 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c7
+ bl_int_51_7 bl_int_50_7 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c8
+ bl_int_51_8 bl_int_50_8 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c9
+ bl_int_51_9 bl_int_50_9 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c10
+ bl_int_51_10 bl_int_50_10 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c11
+ bl_int_51_11 bl_int_50_11 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c12
+ bl_int_51_12 bl_int_50_12 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c13
+ bl_int_51_13 bl_int_50_13 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c14
+ bl_int_51_14 bl_int_50_14 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c15
+ bl_int_51_15 bl_int_50_15 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c16
+ bl_int_51_16 bl_int_50_16 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c17
+ bl_int_51_17 bl_int_50_17 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c18
+ bl_int_51_18 bl_int_50_18 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c19
+ bl_int_51_19 bl_int_50_19 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c20
+ bl_int_51_20 bl_int_50_20 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c21
+ bl_int_51_21 bl_int_50_21 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c22
+ bl_int_51_22 bl_int_50_22 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c23
+ bl_int_51_23 bl_int_50_23 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c24
+ bl_int_51_24 bl_int_50_24 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c25
+ bl_int_51_25 bl_int_50_25 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c26
+ bl_int_51_26 bl_int_50_26 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c27
+ bl_int_51_27 bl_int_50_27 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c28
+ bl_int_51_28 bl_int_50_28 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c29
+ bl_int_51_29 bl_int_50_29 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c30
+ bl_int_51_30 bl_int_50_30 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c31
+ bl_int_51_31 bl_int_50_31 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c32
+ bl_int_51_32 bl_int_50_32 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c33
+ bl_int_51_33 bl_int_50_33 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c34
+ bl_int_51_34 bl_int_50_34 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c35
+ bl_int_51_35 bl_int_50_35 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c36
+ bl_int_51_36 bl_int_50_36 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c37
+ bl_int_51_37 bl_int_50_37 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c38
+ bl_int_51_38 bl_int_50_38 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c39
+ bl_int_51_39 bl_int_50_39 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c40
+ bl_int_51_40 bl_int_50_40 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c41
+ bl_int_51_41 bl_int_50_41 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c42
+ bl_int_51_42 bl_int_50_42 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c43
+ bl_int_51_43 bl_int_50_43 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c44
+ bl_int_51_44 bl_int_50_44 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c45
+ bl_int_51_45 bl_int_50_45 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c46
+ bl_int_51_46 bl_int_50_46 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c47
+ bl_int_51_47 bl_int_50_47 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c48
+ bl_int_51_48 bl_int_50_48 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c49
+ bl_int_51_49 bl_int_50_49 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c50
+ bl_int_51_50 bl_int_50_50 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c51
+ bl_int_51_51 bl_int_50_51 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c52
+ bl_int_51_52 bl_int_50_52 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c53
+ bl_int_51_53 bl_int_50_53 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c54
+ bl_int_51_54 bl_int_50_54 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c55
+ bl_int_51_55 bl_int_50_55 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c56
+ bl_int_51_56 bl_int_50_56 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c57
+ bl_int_51_57 bl_int_50_57 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c58
+ bl_int_51_58 bl_int_50_58 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c59
+ bl_int_51_59 bl_int_50_59 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c60
+ bl_int_51_60 bl_int_50_60 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c61
+ bl_int_51_61 bl_int_50_61 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c62
+ bl_int_51_62 bl_int_50_62 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c63
+ bl_int_51_63 bl_int_50_63 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c64
+ bl_int_51_64 bl_int_50_64 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c65
+ bl_int_51_65 bl_int_50_65 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c66
+ bl_int_51_66 bl_int_50_66 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c67
+ bl_int_51_67 bl_int_50_67 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c68
+ bl_int_51_68 bl_int_50_68 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c69
+ bl_int_51_69 bl_int_50_69 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c70
+ bl_int_51_70 bl_int_50_70 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c71
+ bl_int_51_71 bl_int_50_71 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c72
+ bl_int_51_72 bl_int_50_72 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c73
+ bl_int_51_73 bl_int_50_73 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c74
+ bl_int_51_74 bl_int_50_74 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c75
+ bl_int_51_75 bl_int_50_75 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c76
+ bl_int_51_76 bl_int_50_76 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c77
+ bl_int_51_77 bl_int_50_77 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c78
+ bl_int_51_78 bl_int_50_78 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c79
+ bl_int_51_79 bl_int_50_79 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c80
+ bl_int_51_80 bl_int_50_80 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c81
+ bl_int_51_81 bl_int_50_81 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c82
+ bl_int_51_82 bl_int_50_82 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c83
+ bl_int_51_83 bl_int_50_83 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c84
+ bl_int_51_84 bl_int_50_84 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c85
+ bl_int_51_85 bl_int_50_85 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c86
+ bl_int_51_86 bl_int_50_86 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c87
+ bl_int_51_87 bl_int_50_87 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c88
+ bl_int_51_88 bl_int_50_88 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c89
+ bl_int_51_89 bl_int_50_89 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c90
+ bl_int_51_90 bl_int_50_90 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c91
+ bl_int_51_91 bl_int_50_91 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c92
+ bl_int_51_92 bl_int_50_92 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c93
+ bl_int_51_93 bl_int_50_93 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c94
+ bl_int_51_94 bl_int_50_94 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c95
+ bl_int_51_95 bl_int_50_95 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c96
+ bl_int_51_96 bl_int_50_96 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c97
+ bl_int_51_97 bl_int_50_97 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c98
+ bl_int_51_98 bl_int_50_98 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c99
+ bl_int_51_99 bl_int_50_99 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c100
+ bl_int_51_100 bl_int_50_100 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c101
+ bl_int_51_101 bl_int_50_101 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c102
+ bl_int_51_102 bl_int_50_102 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c103
+ bl_int_51_103 bl_int_50_103 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c104
+ bl_int_51_104 bl_int_50_104 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c105
+ bl_int_51_105 bl_int_50_105 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c106
+ bl_int_51_106 bl_int_50_106 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c107
+ bl_int_51_107 bl_int_50_107 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c108
+ bl_int_51_108 bl_int_50_108 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c109
+ bl_int_51_109 bl_int_50_109 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c110
+ bl_int_51_110 bl_int_50_110 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c111
+ bl_int_51_111 bl_int_50_111 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c112
+ bl_int_51_112 bl_int_50_112 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c113
+ bl_int_51_113 bl_int_50_113 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c114
+ bl_int_51_114 bl_int_50_114 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c115
+ bl_int_51_115 bl_int_50_115 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c116
+ bl_int_51_116 bl_int_50_116 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c117
+ bl_int_51_117 bl_int_50_117 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c118
+ bl_int_51_118 bl_int_50_118 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c119
+ bl_int_51_119 bl_int_50_119 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c120
+ bl_int_51_120 bl_int_50_120 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c121
+ bl_int_51_121 bl_int_50_121 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c122
+ bl_int_51_122 bl_int_50_122 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c123
+ bl_int_51_123 bl_int_50_123 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c124
+ bl_int_51_124 bl_int_50_124 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c125
+ bl_int_51_125 bl_int_50_125 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c126
+ bl_int_51_126 bl_int_50_126 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c127
+ bl_int_51_127 bl_int_50_127 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c128
+ bl_int_51_128 bl_int_50_128 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c129
+ bl_int_51_129 bl_int_50_129 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c130
+ bl_int_51_130 bl_int_50_130 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c131
+ bl_int_51_131 bl_int_50_131 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c132
+ bl_int_51_132 bl_int_50_132 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c133
+ bl_int_51_133 bl_int_50_133 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c134
+ bl_int_51_134 bl_int_50_134 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c135
+ bl_int_51_135 bl_int_50_135 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c136
+ bl_int_51_136 bl_int_50_136 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c137
+ bl_int_51_137 bl_int_50_137 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c138
+ bl_int_51_138 bl_int_50_138 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c139
+ bl_int_51_139 bl_int_50_139 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c140
+ bl_int_51_140 bl_int_50_140 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c141
+ bl_int_51_141 bl_int_50_141 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c142
+ bl_int_51_142 bl_int_50_142 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c143
+ bl_int_51_143 bl_int_50_143 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c144
+ bl_int_51_144 bl_int_50_144 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c145
+ bl_int_51_145 bl_int_50_145 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c146
+ bl_int_51_146 bl_int_50_146 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c147
+ bl_int_51_147 bl_int_50_147 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c148
+ bl_int_51_148 bl_int_50_148 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c149
+ bl_int_51_149 bl_int_50_149 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c150
+ bl_int_51_150 bl_int_50_150 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c151
+ bl_int_51_151 bl_int_50_151 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c152
+ bl_int_51_152 bl_int_50_152 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c153
+ bl_int_51_153 bl_int_50_153 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c154
+ bl_int_51_154 bl_int_50_154 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c155
+ bl_int_51_155 bl_int_50_155 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c156
+ bl_int_51_156 bl_int_50_156 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c157
+ bl_int_51_157 bl_int_50_157 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c158
+ bl_int_51_158 bl_int_50_158 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c159
+ bl_int_51_159 bl_int_50_159 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c160
+ bl_int_51_160 bl_int_50_160 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c161
+ bl_int_51_161 bl_int_50_161 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c162
+ bl_int_51_162 bl_int_50_162 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c163
+ bl_int_51_163 bl_int_50_163 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c164
+ bl_int_51_164 bl_int_50_164 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c165
+ bl_int_51_165 bl_int_50_165 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c166
+ bl_int_51_166 bl_int_50_166 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c167
+ bl_int_51_167 bl_int_50_167 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c168
+ bl_int_51_168 bl_int_50_168 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c169
+ bl_int_51_169 bl_int_50_169 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c170
+ bl_int_51_170 bl_int_50_170 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c171
+ bl_int_51_171 bl_int_50_171 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c172
+ bl_int_51_172 bl_int_50_172 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c173
+ bl_int_51_173 bl_int_50_173 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c174
+ bl_int_51_174 bl_int_50_174 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c175
+ bl_int_51_175 bl_int_50_175 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c176
+ bl_int_51_176 bl_int_50_176 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c177
+ bl_int_51_177 bl_int_50_177 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c178
+ bl_int_51_178 bl_int_50_178 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c179
+ bl_int_51_179 bl_int_50_179 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c180
+ bl_int_51_180 bl_int_50_180 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c181
+ bl_int_51_181 bl_int_50_181 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c182
+ bl_int_51_182 bl_int_50_182 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r51_c183
+ bl_int_51_183 bl_int_50_183 wl_0_51 gnd
+ sram_rom_base_one_cell
Xbit_r52_c0
+ bl_int_52_0 bl_int_51_0 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c1
+ bl_int_52_1 bl_int_51_1 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c2
+ bl_int_52_2 bl_int_51_2 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c3
+ bl_int_52_3 bl_int_51_3 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c4
+ bl_int_52_4 bl_int_51_4 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c5
+ bl_int_52_5 bl_int_51_5 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c6
+ bl_int_52_6 bl_int_51_6 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c7
+ bl_int_52_7 bl_int_51_7 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c8
+ bl_int_52_8 bl_int_51_8 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c9
+ bl_int_52_9 bl_int_51_9 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c10
+ bl_int_52_10 bl_int_51_10 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c11
+ bl_int_52_11 bl_int_51_11 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c12
+ bl_int_52_12 bl_int_51_12 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c13
+ bl_int_52_13 bl_int_51_13 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c14
+ bl_int_52_14 bl_int_51_14 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c15
+ bl_int_52_15 bl_int_51_15 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c16
+ bl_int_52_16 bl_int_51_16 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c17
+ bl_int_52_17 bl_int_51_17 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c18
+ bl_int_52_18 bl_int_51_18 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c19
+ bl_int_52_19 bl_int_51_19 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c20
+ bl_int_52_20 bl_int_51_20 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c21
+ bl_int_52_21 bl_int_51_21 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c22
+ bl_int_52_22 bl_int_51_22 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c23
+ bl_int_52_23 bl_int_51_23 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c24
+ bl_int_52_24 bl_int_51_24 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c25
+ bl_int_52_25 bl_int_51_25 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c26
+ bl_int_52_26 bl_int_51_26 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c27
+ bl_int_52_27 bl_int_51_27 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c28
+ bl_int_52_28 bl_int_51_28 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c29
+ bl_int_52_29 bl_int_51_29 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c30
+ bl_int_52_30 bl_int_51_30 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c31
+ bl_int_52_31 bl_int_51_31 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c32
+ bl_int_52_32 bl_int_51_32 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c33
+ bl_int_52_33 bl_int_51_33 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c34
+ bl_int_52_34 bl_int_51_34 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c35
+ bl_int_52_35 bl_int_51_35 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c36
+ bl_int_52_36 bl_int_51_36 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c37
+ bl_int_52_37 bl_int_51_37 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c38
+ bl_int_52_38 bl_int_51_38 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c39
+ bl_int_52_39 bl_int_51_39 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c40
+ bl_int_52_40 bl_int_51_40 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c41
+ bl_int_52_41 bl_int_51_41 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c42
+ bl_int_52_42 bl_int_51_42 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c43
+ bl_int_52_43 bl_int_51_43 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c44
+ bl_int_52_44 bl_int_51_44 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c45
+ bl_int_52_45 bl_int_51_45 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c46
+ bl_int_52_46 bl_int_51_46 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c47
+ bl_int_52_47 bl_int_51_47 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c48
+ bl_int_52_48 bl_int_51_48 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c49
+ bl_int_52_49 bl_int_51_49 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c50
+ bl_int_52_50 bl_int_51_50 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c51
+ bl_int_52_51 bl_int_51_51 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c52
+ bl_int_52_52 bl_int_51_52 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c53
+ bl_int_52_53 bl_int_51_53 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c54
+ bl_int_52_54 bl_int_51_54 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c55
+ bl_int_52_55 bl_int_51_55 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c56
+ bl_int_52_56 bl_int_51_56 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c57
+ bl_int_52_57 bl_int_51_57 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c58
+ bl_int_52_58 bl_int_51_58 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c59
+ bl_int_52_59 bl_int_51_59 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c60
+ bl_int_52_60 bl_int_51_60 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c61
+ bl_int_52_61 bl_int_51_61 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c62
+ bl_int_52_62 bl_int_51_62 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c63
+ bl_int_52_63 bl_int_51_63 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c64
+ bl_int_52_64 bl_int_51_64 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c65
+ bl_int_52_65 bl_int_51_65 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c66
+ bl_int_52_66 bl_int_51_66 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c67
+ bl_int_52_67 bl_int_51_67 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c68
+ bl_int_52_68 bl_int_51_68 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c69
+ bl_int_52_69 bl_int_51_69 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c70
+ bl_int_52_70 bl_int_51_70 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c71
+ bl_int_52_71 bl_int_51_71 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c72
+ bl_int_52_72 bl_int_51_72 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c73
+ bl_int_52_73 bl_int_51_73 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c74
+ bl_int_52_74 bl_int_51_74 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c75
+ bl_int_52_75 bl_int_51_75 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c76
+ bl_int_52_76 bl_int_51_76 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c77
+ bl_int_52_77 bl_int_51_77 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c78
+ bl_int_52_78 bl_int_51_78 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c79
+ bl_int_52_79 bl_int_51_79 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c80
+ bl_int_52_80 bl_int_51_80 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c81
+ bl_int_52_81 bl_int_51_81 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c82
+ bl_int_52_82 bl_int_51_82 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c83
+ bl_int_52_83 bl_int_51_83 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c84
+ bl_int_52_84 bl_int_51_84 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c85
+ bl_int_52_85 bl_int_51_85 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c86
+ bl_int_52_86 bl_int_51_86 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c87
+ bl_int_52_87 bl_int_51_87 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c88
+ bl_int_52_88 bl_int_51_88 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c89
+ bl_int_52_89 bl_int_51_89 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c90
+ bl_int_52_90 bl_int_51_90 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c91
+ bl_int_52_91 bl_int_51_91 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c92
+ bl_int_52_92 bl_int_51_92 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c93
+ bl_int_52_93 bl_int_51_93 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c94
+ bl_int_52_94 bl_int_51_94 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c95
+ bl_int_52_95 bl_int_51_95 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c96
+ bl_int_52_96 bl_int_51_96 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c97
+ bl_int_52_97 bl_int_51_97 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c98
+ bl_int_52_98 bl_int_51_98 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c99
+ bl_int_52_99 bl_int_51_99 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c100
+ bl_int_52_100 bl_int_51_100 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c101
+ bl_int_52_101 bl_int_51_101 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c102
+ bl_int_52_102 bl_int_51_102 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c103
+ bl_int_52_103 bl_int_51_103 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c104
+ bl_int_52_104 bl_int_51_104 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c105
+ bl_int_52_105 bl_int_51_105 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c106
+ bl_int_52_106 bl_int_51_106 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c107
+ bl_int_52_107 bl_int_51_107 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c108
+ bl_int_52_108 bl_int_51_108 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c109
+ bl_int_52_109 bl_int_51_109 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c110
+ bl_int_52_110 bl_int_51_110 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c111
+ bl_int_52_111 bl_int_51_111 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c112
+ bl_int_52_112 bl_int_51_112 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c113
+ bl_int_52_113 bl_int_51_113 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c114
+ bl_int_52_114 bl_int_51_114 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c115
+ bl_int_52_115 bl_int_51_115 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c116
+ bl_int_52_116 bl_int_51_116 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c117
+ bl_int_52_117 bl_int_51_117 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c118
+ bl_int_52_118 bl_int_51_118 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c119
+ bl_int_52_119 bl_int_51_119 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c120
+ bl_int_52_120 bl_int_51_120 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c121
+ bl_int_52_121 bl_int_51_121 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c122
+ bl_int_52_122 bl_int_51_122 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c123
+ bl_int_52_123 bl_int_51_123 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c124
+ bl_int_52_124 bl_int_51_124 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c125
+ bl_int_52_125 bl_int_51_125 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c126
+ bl_int_52_126 bl_int_51_126 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c127
+ bl_int_52_127 bl_int_51_127 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c128
+ bl_int_52_128 bl_int_51_128 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c129
+ bl_int_52_129 bl_int_51_129 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c130
+ bl_int_52_130 bl_int_51_130 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c131
+ bl_int_52_131 bl_int_51_131 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c132
+ bl_int_52_132 bl_int_51_132 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c133
+ bl_int_52_133 bl_int_51_133 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c134
+ bl_int_52_134 bl_int_51_134 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c135
+ bl_int_52_135 bl_int_51_135 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c136
+ bl_int_52_136 bl_int_51_136 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c137
+ bl_int_52_137 bl_int_51_137 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c138
+ bl_int_52_138 bl_int_51_138 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c139
+ bl_int_52_139 bl_int_51_139 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c140
+ bl_int_52_140 bl_int_51_140 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c141
+ bl_int_52_141 bl_int_51_141 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c142
+ bl_int_52_142 bl_int_51_142 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c143
+ bl_int_52_143 bl_int_51_143 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c144
+ bl_int_52_144 bl_int_51_144 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c145
+ bl_int_52_145 bl_int_51_145 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c146
+ bl_int_52_146 bl_int_51_146 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c147
+ bl_int_52_147 bl_int_51_147 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c148
+ bl_int_52_148 bl_int_51_148 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c149
+ bl_int_52_149 bl_int_51_149 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c150
+ bl_int_52_150 bl_int_51_150 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c151
+ bl_int_52_151 bl_int_51_151 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c152
+ bl_int_52_152 bl_int_51_152 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c153
+ bl_int_52_153 bl_int_51_153 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c154
+ bl_int_52_154 bl_int_51_154 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c155
+ bl_int_52_155 bl_int_51_155 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c156
+ bl_int_52_156 bl_int_51_156 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c157
+ bl_int_52_157 bl_int_51_157 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c158
+ bl_int_52_158 bl_int_51_158 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c159
+ bl_int_52_159 bl_int_51_159 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c160
+ bl_int_52_160 bl_int_51_160 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c161
+ bl_int_52_161 bl_int_51_161 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c162
+ bl_int_52_162 bl_int_51_162 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c163
+ bl_int_52_163 bl_int_51_163 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c164
+ bl_int_52_164 bl_int_51_164 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c165
+ bl_int_52_165 bl_int_51_165 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c166
+ bl_int_52_166 bl_int_51_166 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c167
+ bl_int_52_167 bl_int_51_167 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c168
+ bl_int_52_168 bl_int_51_168 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c169
+ bl_int_52_169 bl_int_51_169 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c170
+ bl_int_52_170 bl_int_51_170 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c171
+ bl_int_52_171 bl_int_51_171 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c172
+ bl_int_52_172 bl_int_51_172 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c173
+ bl_int_52_173 bl_int_51_173 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c174
+ bl_int_52_174 bl_int_51_174 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c175
+ bl_int_52_175 bl_int_51_175 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c176
+ bl_int_52_176 bl_int_51_176 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c177
+ bl_int_52_177 bl_int_51_177 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c178
+ bl_int_52_178 bl_int_51_178 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c179
+ bl_int_52_179 bl_int_51_179 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c180
+ bl_int_52_180 bl_int_51_180 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c181
+ bl_int_52_181 bl_int_51_181 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c182
+ bl_int_52_182 bl_int_51_182 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r52_c183
+ bl_int_52_183 bl_int_51_183 wl_0_52 gnd
+ sram_rom_base_one_cell
Xbit_r53_c0
+ bl_int_53_0 bl_int_52_0 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c1
+ bl_int_53_1 bl_int_52_1 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c2
+ bl_int_53_2 bl_int_52_2 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c3
+ bl_int_53_3 bl_int_52_3 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c4
+ bl_int_53_4 bl_int_52_4 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c5
+ bl_int_53_5 bl_int_52_5 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c6
+ bl_int_53_6 bl_int_52_6 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c7
+ bl_int_53_7 bl_int_52_7 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c8
+ bl_int_53_8 bl_int_52_8 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c9
+ bl_int_53_9 bl_int_52_9 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c10
+ bl_int_53_10 bl_int_52_10 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c11
+ bl_int_53_11 bl_int_52_11 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c12
+ bl_int_53_12 bl_int_52_12 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c13
+ bl_int_53_13 bl_int_52_13 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c14
+ bl_int_53_14 bl_int_52_14 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c15
+ bl_int_53_15 bl_int_52_15 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c16
+ bl_int_53_16 bl_int_52_16 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c17
+ bl_int_53_17 bl_int_52_17 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c18
+ bl_int_53_18 bl_int_52_18 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c19
+ bl_int_53_19 bl_int_52_19 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c20
+ bl_int_53_20 bl_int_52_20 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c21
+ bl_int_53_21 bl_int_52_21 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c22
+ bl_int_53_22 bl_int_52_22 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c23
+ bl_int_53_23 bl_int_52_23 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c24
+ bl_int_53_24 bl_int_52_24 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c25
+ bl_int_53_25 bl_int_52_25 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c26
+ bl_int_53_26 bl_int_52_26 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c27
+ bl_int_53_27 bl_int_52_27 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c28
+ bl_int_53_28 bl_int_52_28 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c29
+ bl_int_53_29 bl_int_52_29 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c30
+ bl_int_53_30 bl_int_52_30 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c31
+ bl_int_53_31 bl_int_52_31 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c32
+ bl_int_53_32 bl_int_52_32 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c33
+ bl_int_53_33 bl_int_52_33 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c34
+ bl_int_53_34 bl_int_52_34 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c35
+ bl_int_53_35 bl_int_52_35 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c36
+ bl_int_53_36 bl_int_52_36 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c37
+ bl_int_53_37 bl_int_52_37 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c38
+ bl_int_53_38 bl_int_52_38 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c39
+ bl_int_53_39 bl_int_52_39 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c40
+ bl_int_53_40 bl_int_52_40 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c41
+ bl_int_53_41 bl_int_52_41 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c42
+ bl_int_53_42 bl_int_52_42 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c43
+ bl_int_53_43 bl_int_52_43 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c44
+ bl_int_53_44 bl_int_52_44 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c45
+ bl_int_53_45 bl_int_52_45 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c46
+ bl_int_53_46 bl_int_52_46 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c47
+ bl_int_53_47 bl_int_52_47 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c48
+ bl_int_53_48 bl_int_52_48 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c49
+ bl_int_53_49 bl_int_52_49 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c50
+ bl_int_53_50 bl_int_52_50 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c51
+ bl_int_53_51 bl_int_52_51 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c52
+ bl_int_53_52 bl_int_52_52 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c53
+ bl_int_53_53 bl_int_52_53 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c54
+ bl_int_53_54 bl_int_52_54 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c55
+ bl_int_53_55 bl_int_52_55 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c56
+ bl_int_53_56 bl_int_52_56 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c57
+ bl_int_53_57 bl_int_52_57 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c58
+ bl_int_53_58 bl_int_52_58 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c59
+ bl_int_53_59 bl_int_52_59 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c60
+ bl_int_53_60 bl_int_52_60 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c61
+ bl_int_53_61 bl_int_52_61 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c62
+ bl_int_53_62 bl_int_52_62 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c63
+ bl_int_53_63 bl_int_52_63 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c64
+ bl_int_53_64 bl_int_52_64 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c65
+ bl_int_53_65 bl_int_52_65 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c66
+ bl_int_53_66 bl_int_52_66 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c67
+ bl_int_53_67 bl_int_52_67 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c68
+ bl_int_53_68 bl_int_52_68 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c69
+ bl_int_53_69 bl_int_52_69 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c70
+ bl_int_53_70 bl_int_52_70 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c71
+ bl_int_53_71 bl_int_52_71 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c72
+ bl_int_53_72 bl_int_52_72 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c73
+ bl_int_53_73 bl_int_52_73 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c74
+ bl_int_53_74 bl_int_52_74 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c75
+ bl_int_53_75 bl_int_52_75 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c76
+ bl_int_53_76 bl_int_52_76 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c77
+ bl_int_53_77 bl_int_52_77 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c78
+ bl_int_53_78 bl_int_52_78 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c79
+ bl_int_53_79 bl_int_52_79 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c80
+ bl_int_53_80 bl_int_52_80 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c81
+ bl_int_53_81 bl_int_52_81 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c82
+ bl_int_53_82 bl_int_52_82 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c83
+ bl_int_53_83 bl_int_52_83 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c84
+ bl_int_53_84 bl_int_52_84 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c85
+ bl_int_53_85 bl_int_52_85 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c86
+ bl_int_53_86 bl_int_52_86 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c87
+ bl_int_53_87 bl_int_52_87 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c88
+ bl_int_53_88 bl_int_52_88 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c89
+ bl_int_53_89 bl_int_52_89 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c90
+ bl_int_53_90 bl_int_52_90 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c91
+ bl_int_53_91 bl_int_52_91 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c92
+ bl_int_53_92 bl_int_52_92 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c93
+ bl_int_53_93 bl_int_52_93 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c94
+ bl_int_53_94 bl_int_52_94 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c95
+ bl_int_53_95 bl_int_52_95 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c96
+ bl_int_53_96 bl_int_52_96 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c97
+ bl_int_53_97 bl_int_52_97 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c98
+ bl_int_53_98 bl_int_52_98 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c99
+ bl_int_53_99 bl_int_52_99 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c100
+ bl_int_53_100 bl_int_52_100 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c101
+ bl_int_53_101 bl_int_52_101 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c102
+ bl_int_53_102 bl_int_52_102 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c103
+ bl_int_53_103 bl_int_52_103 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c104
+ bl_int_53_104 bl_int_52_104 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c105
+ bl_int_53_105 bl_int_52_105 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c106
+ bl_int_53_106 bl_int_52_106 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c107
+ bl_int_53_107 bl_int_52_107 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c108
+ bl_int_53_108 bl_int_52_108 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c109
+ bl_int_53_109 bl_int_52_109 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c110
+ bl_int_53_110 bl_int_52_110 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c111
+ bl_int_53_111 bl_int_52_111 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c112
+ bl_int_53_112 bl_int_52_112 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c113
+ bl_int_53_113 bl_int_52_113 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c114
+ bl_int_53_114 bl_int_52_114 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c115
+ bl_int_53_115 bl_int_52_115 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c116
+ bl_int_53_116 bl_int_52_116 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c117
+ bl_int_53_117 bl_int_52_117 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c118
+ bl_int_53_118 bl_int_52_118 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c119
+ bl_int_53_119 bl_int_52_119 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c120
+ bl_int_53_120 bl_int_52_120 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c121
+ bl_int_53_121 bl_int_52_121 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c122
+ bl_int_53_122 bl_int_52_122 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c123
+ bl_int_53_123 bl_int_52_123 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c124
+ bl_int_53_124 bl_int_52_124 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c125
+ bl_int_53_125 bl_int_52_125 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c126
+ bl_int_53_126 bl_int_52_126 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c127
+ bl_int_53_127 bl_int_52_127 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c128
+ bl_int_53_128 bl_int_52_128 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c129
+ bl_int_53_129 bl_int_52_129 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c130
+ bl_int_53_130 bl_int_52_130 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c131
+ bl_int_53_131 bl_int_52_131 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c132
+ bl_int_53_132 bl_int_52_132 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c133
+ bl_int_53_133 bl_int_52_133 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c134
+ bl_int_53_134 bl_int_52_134 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c135
+ bl_int_53_135 bl_int_52_135 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c136
+ bl_int_53_136 bl_int_52_136 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c137
+ bl_int_53_137 bl_int_52_137 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c138
+ bl_int_53_138 bl_int_52_138 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c139
+ bl_int_53_139 bl_int_52_139 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c140
+ bl_int_53_140 bl_int_52_140 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c141
+ bl_int_53_141 bl_int_52_141 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c142
+ bl_int_53_142 bl_int_52_142 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c143
+ bl_int_53_143 bl_int_52_143 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c144
+ bl_int_53_144 bl_int_52_144 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c145
+ bl_int_53_145 bl_int_52_145 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c146
+ bl_int_53_146 bl_int_52_146 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c147
+ bl_int_53_147 bl_int_52_147 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c148
+ bl_int_53_148 bl_int_52_148 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c149
+ bl_int_53_149 bl_int_52_149 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c150
+ bl_int_53_150 bl_int_52_150 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c151
+ bl_int_53_151 bl_int_52_151 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c152
+ bl_int_53_152 bl_int_52_152 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c153
+ bl_int_53_153 bl_int_52_153 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c154
+ bl_int_53_154 bl_int_52_154 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c155
+ bl_int_53_155 bl_int_52_155 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c156
+ bl_int_53_156 bl_int_52_156 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c157
+ bl_int_53_157 bl_int_52_157 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c158
+ bl_int_53_158 bl_int_52_158 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c159
+ bl_int_53_159 bl_int_52_159 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c160
+ bl_int_53_160 bl_int_52_160 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c161
+ bl_int_53_161 bl_int_52_161 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c162
+ bl_int_53_162 bl_int_52_162 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c163
+ bl_int_53_163 bl_int_52_163 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c164
+ bl_int_53_164 bl_int_52_164 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c165
+ bl_int_53_165 bl_int_52_165 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c166
+ bl_int_53_166 bl_int_52_166 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c167
+ bl_int_53_167 bl_int_52_167 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c168
+ bl_int_53_168 bl_int_52_168 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c169
+ bl_int_53_169 bl_int_52_169 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c170
+ bl_int_53_170 bl_int_52_170 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c171
+ bl_int_53_171 bl_int_52_171 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c172
+ bl_int_53_172 bl_int_52_172 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c173
+ bl_int_53_173 bl_int_52_173 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c174
+ bl_int_53_174 bl_int_52_174 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c175
+ bl_int_53_175 bl_int_52_175 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c176
+ bl_int_53_176 bl_int_52_176 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c177
+ bl_int_53_177 bl_int_52_177 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c178
+ bl_int_53_178 bl_int_52_178 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c179
+ bl_int_53_179 bl_int_52_179 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c180
+ bl_int_53_180 bl_int_52_180 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c181
+ bl_int_53_181 bl_int_52_181 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c182
+ bl_int_53_182 bl_int_52_182 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r53_c183
+ bl_int_53_183 bl_int_52_183 wl_0_53 gnd
+ sram_rom_base_one_cell
Xbit_r54_c0
+ bl_int_54_0 bl_int_53_0 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c1
+ bl_int_54_1 bl_int_53_1 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c2
+ bl_int_54_2 bl_int_53_2 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c3
+ bl_int_54_3 bl_int_53_3 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c4
+ bl_int_54_4 bl_int_53_4 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c5
+ bl_int_54_5 bl_int_53_5 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c6
+ bl_int_54_6 bl_int_53_6 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c7
+ bl_int_54_7 bl_int_53_7 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c8
+ bl_int_54_8 bl_int_53_8 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c9
+ bl_int_54_9 bl_int_53_9 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c10
+ bl_int_54_10 bl_int_53_10 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c11
+ bl_int_54_11 bl_int_53_11 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c12
+ bl_int_54_12 bl_int_53_12 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c13
+ bl_int_54_13 bl_int_53_13 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c14
+ bl_int_54_14 bl_int_53_14 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c15
+ bl_int_54_15 bl_int_53_15 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c16
+ bl_int_54_16 bl_int_53_16 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c17
+ bl_int_54_17 bl_int_53_17 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c18
+ bl_int_54_18 bl_int_53_18 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c19
+ bl_int_54_19 bl_int_53_19 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c20
+ bl_int_54_20 bl_int_53_20 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c21
+ bl_int_54_21 bl_int_53_21 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c22
+ bl_int_54_22 bl_int_53_22 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c23
+ bl_int_54_23 bl_int_53_23 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c24
+ bl_int_54_24 bl_int_53_24 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c25
+ bl_int_54_25 bl_int_53_25 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c26
+ bl_int_54_26 bl_int_53_26 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c27
+ bl_int_54_27 bl_int_53_27 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c28
+ bl_int_54_28 bl_int_53_28 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c29
+ bl_int_54_29 bl_int_53_29 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c30
+ bl_int_54_30 bl_int_53_30 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c31
+ bl_int_54_31 bl_int_53_31 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c32
+ bl_int_54_32 bl_int_53_32 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c33
+ bl_int_54_33 bl_int_53_33 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c34
+ bl_int_54_34 bl_int_53_34 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c35
+ bl_int_54_35 bl_int_53_35 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c36
+ bl_int_54_36 bl_int_53_36 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c37
+ bl_int_54_37 bl_int_53_37 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c38
+ bl_int_54_38 bl_int_53_38 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c39
+ bl_int_54_39 bl_int_53_39 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c40
+ bl_int_54_40 bl_int_53_40 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c41
+ bl_int_54_41 bl_int_53_41 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c42
+ bl_int_54_42 bl_int_53_42 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c43
+ bl_int_54_43 bl_int_53_43 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c44
+ bl_int_54_44 bl_int_53_44 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c45
+ bl_int_54_45 bl_int_53_45 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c46
+ bl_int_54_46 bl_int_53_46 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c47
+ bl_int_54_47 bl_int_53_47 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c48
+ bl_int_54_48 bl_int_53_48 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c49
+ bl_int_54_49 bl_int_53_49 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c50
+ bl_int_54_50 bl_int_53_50 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c51
+ bl_int_54_51 bl_int_53_51 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c52
+ bl_int_54_52 bl_int_53_52 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c53
+ bl_int_54_53 bl_int_53_53 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c54
+ bl_int_54_54 bl_int_53_54 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c55
+ bl_int_54_55 bl_int_53_55 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c56
+ bl_int_54_56 bl_int_53_56 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c57
+ bl_int_54_57 bl_int_53_57 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c58
+ bl_int_54_58 bl_int_53_58 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c59
+ bl_int_54_59 bl_int_53_59 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c60
+ bl_int_54_60 bl_int_53_60 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c61
+ bl_int_54_61 bl_int_53_61 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c62
+ bl_int_54_62 bl_int_53_62 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c63
+ bl_int_54_63 bl_int_53_63 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c64
+ bl_int_54_64 bl_int_53_64 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c65
+ bl_int_54_65 bl_int_53_65 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c66
+ bl_int_54_66 bl_int_53_66 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c67
+ bl_int_54_67 bl_int_53_67 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c68
+ bl_int_54_68 bl_int_53_68 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c69
+ bl_int_54_69 bl_int_53_69 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c70
+ bl_int_54_70 bl_int_53_70 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c71
+ bl_int_54_71 bl_int_53_71 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c72
+ bl_int_54_72 bl_int_53_72 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c73
+ bl_int_54_73 bl_int_53_73 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c74
+ bl_int_54_74 bl_int_53_74 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c75
+ bl_int_54_75 bl_int_53_75 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c76
+ bl_int_54_76 bl_int_53_76 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c77
+ bl_int_54_77 bl_int_53_77 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c78
+ bl_int_54_78 bl_int_53_78 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c79
+ bl_int_54_79 bl_int_53_79 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c80
+ bl_int_54_80 bl_int_53_80 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c81
+ bl_int_54_81 bl_int_53_81 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c82
+ bl_int_54_82 bl_int_53_82 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c83
+ bl_int_54_83 bl_int_53_83 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c84
+ bl_int_54_84 bl_int_53_84 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c85
+ bl_int_54_85 bl_int_53_85 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c86
+ bl_int_54_86 bl_int_53_86 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c87
+ bl_int_54_87 bl_int_53_87 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c88
+ bl_int_54_88 bl_int_53_88 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c89
+ bl_int_54_89 bl_int_53_89 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c90
+ bl_int_54_90 bl_int_53_90 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c91
+ bl_int_54_91 bl_int_53_91 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c92
+ bl_int_54_92 bl_int_53_92 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c93
+ bl_int_54_93 bl_int_53_93 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c94
+ bl_int_54_94 bl_int_53_94 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c95
+ bl_int_54_95 bl_int_53_95 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c96
+ bl_int_54_96 bl_int_53_96 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c97
+ bl_int_54_97 bl_int_53_97 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c98
+ bl_int_54_98 bl_int_53_98 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c99
+ bl_int_54_99 bl_int_53_99 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c100
+ bl_int_54_100 bl_int_53_100 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c101
+ bl_int_54_101 bl_int_53_101 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c102
+ bl_int_54_102 bl_int_53_102 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c103
+ bl_int_54_103 bl_int_53_103 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c104
+ bl_int_54_104 bl_int_53_104 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c105
+ bl_int_54_105 bl_int_53_105 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c106
+ bl_int_54_106 bl_int_53_106 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c107
+ bl_int_54_107 bl_int_53_107 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c108
+ bl_int_54_108 bl_int_53_108 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c109
+ bl_int_54_109 bl_int_53_109 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c110
+ bl_int_54_110 bl_int_53_110 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c111
+ bl_int_54_111 bl_int_53_111 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c112
+ bl_int_54_112 bl_int_53_112 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c113
+ bl_int_54_113 bl_int_53_113 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c114
+ bl_int_54_114 bl_int_53_114 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c115
+ bl_int_54_115 bl_int_53_115 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c116
+ bl_int_54_116 bl_int_53_116 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c117
+ bl_int_54_117 bl_int_53_117 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c118
+ bl_int_54_118 bl_int_53_118 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c119
+ bl_int_54_119 bl_int_53_119 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c120
+ bl_int_54_120 bl_int_53_120 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c121
+ bl_int_54_121 bl_int_53_121 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c122
+ bl_int_54_122 bl_int_53_122 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c123
+ bl_int_54_123 bl_int_53_123 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c124
+ bl_int_54_124 bl_int_53_124 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c125
+ bl_int_54_125 bl_int_53_125 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c126
+ bl_int_54_126 bl_int_53_126 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c127
+ bl_int_54_127 bl_int_53_127 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c128
+ bl_int_54_128 bl_int_53_128 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c129
+ bl_int_54_129 bl_int_53_129 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c130
+ bl_int_54_130 bl_int_53_130 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c131
+ bl_int_54_131 bl_int_53_131 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c132
+ bl_int_54_132 bl_int_53_132 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c133
+ bl_int_54_133 bl_int_53_133 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c134
+ bl_int_54_134 bl_int_53_134 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c135
+ bl_int_54_135 bl_int_53_135 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c136
+ bl_int_54_136 bl_int_53_136 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c137
+ bl_int_54_137 bl_int_53_137 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c138
+ bl_int_54_138 bl_int_53_138 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c139
+ bl_int_54_139 bl_int_53_139 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c140
+ bl_int_54_140 bl_int_53_140 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c141
+ bl_int_54_141 bl_int_53_141 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c142
+ bl_int_54_142 bl_int_53_142 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c143
+ bl_int_54_143 bl_int_53_143 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c144
+ bl_int_54_144 bl_int_53_144 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c145
+ bl_int_54_145 bl_int_53_145 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c146
+ bl_int_54_146 bl_int_53_146 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c147
+ bl_int_54_147 bl_int_53_147 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c148
+ bl_int_54_148 bl_int_53_148 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c149
+ bl_int_54_149 bl_int_53_149 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c150
+ bl_int_54_150 bl_int_53_150 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c151
+ bl_int_54_151 bl_int_53_151 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c152
+ bl_int_54_152 bl_int_53_152 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c153
+ bl_int_54_153 bl_int_53_153 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c154
+ bl_int_54_154 bl_int_53_154 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c155
+ bl_int_54_155 bl_int_53_155 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c156
+ bl_int_54_156 bl_int_53_156 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c157
+ bl_int_54_157 bl_int_53_157 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c158
+ bl_int_54_158 bl_int_53_158 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c159
+ bl_int_54_159 bl_int_53_159 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c160
+ bl_int_54_160 bl_int_53_160 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c161
+ bl_int_54_161 bl_int_53_161 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c162
+ bl_int_54_162 bl_int_53_162 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c163
+ bl_int_54_163 bl_int_53_163 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c164
+ bl_int_54_164 bl_int_53_164 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c165
+ bl_int_54_165 bl_int_53_165 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c166
+ bl_int_54_166 bl_int_53_166 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c167
+ bl_int_54_167 bl_int_53_167 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c168
+ bl_int_54_168 bl_int_53_168 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c169
+ bl_int_54_169 bl_int_53_169 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c170
+ bl_int_54_170 bl_int_53_170 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c171
+ bl_int_54_171 bl_int_53_171 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c172
+ bl_int_54_172 bl_int_53_172 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c173
+ bl_int_54_173 bl_int_53_173 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c174
+ bl_int_54_174 bl_int_53_174 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c175
+ bl_int_54_175 bl_int_53_175 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c176
+ bl_int_54_176 bl_int_53_176 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c177
+ bl_int_54_177 bl_int_53_177 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c178
+ bl_int_54_178 bl_int_53_178 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c179
+ bl_int_54_179 bl_int_53_179 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c180
+ bl_int_54_180 bl_int_53_180 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c181
+ bl_int_54_181 bl_int_53_181 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c182
+ bl_int_54_182 bl_int_53_182 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r54_c183
+ bl_int_54_183 bl_int_53_183 wl_0_54 gnd
+ sram_rom_base_one_cell
Xbit_r55_c0
+ bl_int_55_0 bl_int_54_0 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c1
+ bl_int_55_1 bl_int_54_1 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c2
+ bl_int_55_2 bl_int_54_2 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c3
+ bl_int_55_3 bl_int_54_3 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c4
+ bl_int_55_4 bl_int_54_4 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c5
+ bl_int_55_5 bl_int_54_5 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c6
+ bl_int_55_6 bl_int_54_6 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c7
+ bl_int_55_7 bl_int_54_7 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c8
+ bl_int_55_8 bl_int_54_8 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c9
+ bl_int_55_9 bl_int_54_9 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c10
+ bl_int_55_10 bl_int_54_10 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c11
+ bl_int_55_11 bl_int_54_11 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c12
+ bl_int_55_12 bl_int_54_12 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c13
+ bl_int_55_13 bl_int_54_13 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c14
+ bl_int_55_14 bl_int_54_14 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c15
+ bl_int_55_15 bl_int_54_15 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c16
+ bl_int_55_16 bl_int_54_16 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c17
+ bl_int_55_17 bl_int_54_17 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c18
+ bl_int_55_18 bl_int_54_18 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c19
+ bl_int_55_19 bl_int_54_19 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c20
+ bl_int_55_20 bl_int_54_20 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c21
+ bl_int_55_21 bl_int_54_21 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c22
+ bl_int_55_22 bl_int_54_22 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c23
+ bl_int_55_23 bl_int_54_23 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c24
+ bl_int_55_24 bl_int_54_24 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c25
+ bl_int_55_25 bl_int_54_25 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c26
+ bl_int_55_26 bl_int_54_26 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c27
+ bl_int_55_27 bl_int_54_27 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c28
+ bl_int_55_28 bl_int_54_28 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c29
+ bl_int_55_29 bl_int_54_29 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c30
+ bl_int_55_30 bl_int_54_30 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c31
+ bl_int_55_31 bl_int_54_31 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c32
+ bl_int_55_32 bl_int_54_32 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c33
+ bl_int_55_33 bl_int_54_33 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c34
+ bl_int_55_34 bl_int_54_34 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c35
+ bl_int_55_35 bl_int_54_35 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c36
+ bl_int_55_36 bl_int_54_36 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c37
+ bl_int_55_37 bl_int_54_37 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c38
+ bl_int_55_38 bl_int_54_38 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c39
+ bl_int_55_39 bl_int_54_39 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c40
+ bl_int_55_40 bl_int_54_40 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c41
+ bl_int_55_41 bl_int_54_41 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c42
+ bl_int_55_42 bl_int_54_42 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c43
+ bl_int_55_43 bl_int_54_43 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c44
+ bl_int_55_44 bl_int_54_44 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c45
+ bl_int_55_45 bl_int_54_45 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c46
+ bl_int_55_46 bl_int_54_46 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c47
+ bl_int_55_47 bl_int_54_47 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c48
+ bl_int_55_48 bl_int_54_48 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c49
+ bl_int_55_49 bl_int_54_49 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c50
+ bl_int_55_50 bl_int_54_50 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c51
+ bl_int_55_51 bl_int_54_51 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c52
+ bl_int_55_52 bl_int_54_52 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c53
+ bl_int_55_53 bl_int_54_53 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c54
+ bl_int_55_54 bl_int_54_54 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c55
+ bl_int_55_55 bl_int_54_55 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c56
+ bl_int_55_56 bl_int_54_56 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c57
+ bl_int_55_57 bl_int_54_57 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c58
+ bl_int_55_58 bl_int_54_58 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c59
+ bl_int_55_59 bl_int_54_59 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c60
+ bl_int_55_60 bl_int_54_60 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c61
+ bl_int_55_61 bl_int_54_61 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c62
+ bl_int_55_62 bl_int_54_62 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c63
+ bl_int_55_63 bl_int_54_63 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c64
+ bl_int_55_64 bl_int_54_64 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c65
+ bl_int_55_65 bl_int_54_65 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c66
+ bl_int_55_66 bl_int_54_66 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c67
+ bl_int_55_67 bl_int_54_67 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c68
+ bl_int_55_68 bl_int_54_68 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c69
+ bl_int_55_69 bl_int_54_69 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c70
+ bl_int_55_70 bl_int_54_70 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c71
+ bl_int_55_71 bl_int_54_71 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c72
+ bl_int_55_72 bl_int_54_72 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c73
+ bl_int_55_73 bl_int_54_73 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c74
+ bl_int_55_74 bl_int_54_74 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c75
+ bl_int_55_75 bl_int_54_75 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c76
+ bl_int_55_76 bl_int_54_76 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c77
+ bl_int_55_77 bl_int_54_77 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c78
+ bl_int_55_78 bl_int_54_78 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c79
+ bl_int_55_79 bl_int_54_79 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c80
+ bl_int_55_80 bl_int_54_80 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c81
+ bl_int_55_81 bl_int_54_81 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c82
+ bl_int_55_82 bl_int_54_82 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c83
+ bl_int_55_83 bl_int_54_83 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c84
+ bl_int_55_84 bl_int_54_84 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c85
+ bl_int_55_85 bl_int_54_85 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c86
+ bl_int_55_86 bl_int_54_86 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c87
+ bl_int_55_87 bl_int_54_87 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c88
+ bl_int_55_88 bl_int_54_88 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c89
+ bl_int_55_89 bl_int_54_89 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c90
+ bl_int_55_90 bl_int_54_90 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c91
+ bl_int_55_91 bl_int_54_91 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c92
+ bl_int_55_92 bl_int_54_92 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c93
+ bl_int_55_93 bl_int_54_93 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c94
+ bl_int_55_94 bl_int_54_94 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c95
+ bl_int_55_95 bl_int_54_95 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c96
+ bl_int_55_96 bl_int_54_96 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c97
+ bl_int_55_97 bl_int_54_97 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c98
+ bl_int_55_98 bl_int_54_98 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c99
+ bl_int_55_99 bl_int_54_99 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c100
+ bl_int_55_100 bl_int_54_100 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c101
+ bl_int_55_101 bl_int_54_101 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c102
+ bl_int_55_102 bl_int_54_102 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c103
+ bl_int_55_103 bl_int_54_103 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c104
+ bl_int_55_104 bl_int_54_104 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c105
+ bl_int_55_105 bl_int_54_105 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c106
+ bl_int_55_106 bl_int_54_106 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c107
+ bl_int_55_107 bl_int_54_107 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c108
+ bl_int_55_108 bl_int_54_108 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c109
+ bl_int_55_109 bl_int_54_109 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c110
+ bl_int_55_110 bl_int_54_110 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c111
+ bl_int_55_111 bl_int_54_111 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c112
+ bl_int_55_112 bl_int_54_112 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c113
+ bl_int_55_113 bl_int_54_113 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c114
+ bl_int_55_114 bl_int_54_114 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c115
+ bl_int_55_115 bl_int_54_115 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c116
+ bl_int_55_116 bl_int_54_116 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c117
+ bl_int_55_117 bl_int_54_117 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c118
+ bl_int_55_118 bl_int_54_118 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c119
+ bl_int_55_119 bl_int_54_119 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c120
+ bl_int_55_120 bl_int_54_120 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c121
+ bl_int_55_121 bl_int_54_121 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c122
+ bl_int_55_122 bl_int_54_122 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c123
+ bl_int_55_123 bl_int_54_123 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c124
+ bl_int_55_124 bl_int_54_124 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c125
+ bl_int_55_125 bl_int_54_125 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c126
+ bl_int_55_126 bl_int_54_126 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c127
+ bl_int_55_127 bl_int_54_127 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c128
+ bl_int_55_128 bl_int_54_128 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c129
+ bl_int_55_129 bl_int_54_129 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c130
+ bl_int_55_130 bl_int_54_130 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c131
+ bl_int_55_131 bl_int_54_131 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c132
+ bl_int_55_132 bl_int_54_132 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c133
+ bl_int_55_133 bl_int_54_133 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c134
+ bl_int_55_134 bl_int_54_134 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c135
+ bl_int_55_135 bl_int_54_135 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c136
+ bl_int_55_136 bl_int_54_136 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c137
+ bl_int_55_137 bl_int_54_137 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c138
+ bl_int_55_138 bl_int_54_138 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c139
+ bl_int_55_139 bl_int_54_139 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c140
+ bl_int_55_140 bl_int_54_140 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c141
+ bl_int_55_141 bl_int_54_141 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c142
+ bl_int_55_142 bl_int_54_142 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c143
+ bl_int_55_143 bl_int_54_143 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c144
+ bl_int_55_144 bl_int_54_144 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c145
+ bl_int_55_145 bl_int_54_145 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c146
+ bl_int_55_146 bl_int_54_146 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c147
+ bl_int_55_147 bl_int_54_147 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c148
+ bl_int_55_148 bl_int_54_148 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c149
+ bl_int_55_149 bl_int_54_149 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c150
+ bl_int_55_150 bl_int_54_150 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c151
+ bl_int_55_151 bl_int_54_151 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c152
+ bl_int_55_152 bl_int_54_152 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c153
+ bl_int_55_153 bl_int_54_153 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c154
+ bl_int_55_154 bl_int_54_154 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c155
+ bl_int_55_155 bl_int_54_155 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c156
+ bl_int_55_156 bl_int_54_156 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c157
+ bl_int_55_157 bl_int_54_157 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c158
+ bl_int_55_158 bl_int_54_158 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c159
+ bl_int_55_159 bl_int_54_159 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c160
+ bl_int_55_160 bl_int_54_160 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c161
+ bl_int_55_161 bl_int_54_161 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c162
+ bl_int_55_162 bl_int_54_162 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c163
+ bl_int_55_163 bl_int_54_163 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c164
+ bl_int_55_164 bl_int_54_164 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c165
+ bl_int_55_165 bl_int_54_165 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c166
+ bl_int_55_166 bl_int_54_166 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c167
+ bl_int_55_167 bl_int_54_167 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c168
+ bl_int_55_168 bl_int_54_168 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c169
+ bl_int_55_169 bl_int_54_169 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c170
+ bl_int_55_170 bl_int_54_170 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c171
+ bl_int_55_171 bl_int_54_171 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c172
+ bl_int_55_172 bl_int_54_172 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c173
+ bl_int_55_173 bl_int_54_173 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c174
+ bl_int_55_174 bl_int_54_174 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c175
+ bl_int_55_175 bl_int_54_175 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c176
+ bl_int_55_176 bl_int_54_176 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c177
+ bl_int_55_177 bl_int_54_177 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c178
+ bl_int_55_178 bl_int_54_178 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c179
+ bl_int_55_179 bl_int_54_179 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c180
+ bl_int_55_180 bl_int_54_180 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c181
+ bl_int_55_181 bl_int_54_181 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c182
+ bl_int_55_182 bl_int_54_182 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r55_c183
+ bl_int_55_183 bl_int_54_183 wl_0_55 gnd
+ sram_rom_base_one_cell
Xbit_r56_c0
+ bl_int_56_0 bl_int_55_0 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c1
+ bl_int_56_1 bl_int_55_1 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c2
+ bl_int_56_2 bl_int_55_2 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c3
+ bl_int_56_3 bl_int_55_3 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c4
+ bl_int_56_4 bl_int_55_4 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c5
+ bl_int_56_5 bl_int_55_5 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c6
+ bl_int_56_6 bl_int_55_6 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c7
+ bl_int_56_7 bl_int_55_7 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c8
+ bl_int_56_8 bl_int_55_8 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c9
+ bl_int_56_9 bl_int_55_9 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c10
+ bl_int_56_10 bl_int_55_10 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c11
+ bl_int_56_11 bl_int_55_11 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c12
+ bl_int_56_12 bl_int_55_12 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c13
+ bl_int_56_13 bl_int_55_13 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c14
+ bl_int_56_14 bl_int_55_14 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c15
+ bl_int_56_15 bl_int_55_15 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c16
+ bl_int_56_16 bl_int_55_16 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c17
+ bl_int_56_17 bl_int_55_17 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c18
+ bl_int_56_18 bl_int_55_18 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c19
+ bl_int_56_19 bl_int_55_19 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c20
+ bl_int_56_20 bl_int_55_20 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c21
+ bl_int_56_21 bl_int_55_21 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c22
+ bl_int_56_22 bl_int_55_22 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c23
+ bl_int_56_23 bl_int_55_23 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c24
+ bl_int_56_24 bl_int_55_24 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c25
+ bl_int_56_25 bl_int_55_25 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c26
+ bl_int_56_26 bl_int_55_26 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c27
+ bl_int_56_27 bl_int_55_27 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c28
+ bl_int_56_28 bl_int_55_28 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c29
+ bl_int_56_29 bl_int_55_29 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c30
+ bl_int_56_30 bl_int_55_30 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c31
+ bl_int_56_31 bl_int_55_31 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c32
+ bl_int_56_32 bl_int_55_32 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c33
+ bl_int_56_33 bl_int_55_33 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c34
+ bl_int_56_34 bl_int_55_34 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c35
+ bl_int_56_35 bl_int_55_35 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c36
+ bl_int_56_36 bl_int_55_36 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c37
+ bl_int_56_37 bl_int_55_37 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c38
+ bl_int_56_38 bl_int_55_38 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c39
+ bl_int_56_39 bl_int_55_39 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c40
+ bl_int_56_40 bl_int_55_40 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c41
+ bl_int_56_41 bl_int_55_41 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c42
+ bl_int_56_42 bl_int_55_42 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c43
+ bl_int_56_43 bl_int_55_43 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c44
+ bl_int_56_44 bl_int_55_44 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c45
+ bl_int_56_45 bl_int_55_45 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c46
+ bl_int_56_46 bl_int_55_46 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c47
+ bl_int_56_47 bl_int_55_47 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c48
+ bl_int_56_48 bl_int_55_48 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c49
+ bl_int_56_49 bl_int_55_49 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c50
+ bl_int_56_50 bl_int_55_50 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c51
+ bl_int_56_51 bl_int_55_51 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c52
+ bl_int_56_52 bl_int_55_52 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c53
+ bl_int_56_53 bl_int_55_53 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c54
+ bl_int_56_54 bl_int_55_54 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c55
+ bl_int_56_55 bl_int_55_55 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c56
+ bl_int_56_56 bl_int_55_56 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c57
+ bl_int_56_57 bl_int_55_57 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c58
+ bl_int_56_58 bl_int_55_58 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c59
+ bl_int_56_59 bl_int_55_59 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c60
+ bl_int_56_60 bl_int_55_60 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c61
+ bl_int_56_61 bl_int_55_61 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c62
+ bl_int_56_62 bl_int_55_62 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c63
+ bl_int_56_63 bl_int_55_63 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c64
+ bl_int_56_64 bl_int_55_64 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c65
+ bl_int_56_65 bl_int_55_65 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c66
+ bl_int_56_66 bl_int_55_66 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c67
+ bl_int_56_67 bl_int_55_67 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c68
+ bl_int_56_68 bl_int_55_68 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c69
+ bl_int_56_69 bl_int_55_69 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c70
+ bl_int_56_70 bl_int_55_70 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c71
+ bl_int_56_71 bl_int_55_71 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c72
+ bl_int_56_72 bl_int_55_72 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c73
+ bl_int_56_73 bl_int_55_73 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c74
+ bl_int_56_74 bl_int_55_74 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c75
+ bl_int_56_75 bl_int_55_75 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c76
+ bl_int_56_76 bl_int_55_76 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c77
+ bl_int_56_77 bl_int_55_77 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c78
+ bl_int_56_78 bl_int_55_78 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c79
+ bl_int_56_79 bl_int_55_79 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c80
+ bl_int_56_80 bl_int_55_80 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c81
+ bl_int_56_81 bl_int_55_81 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c82
+ bl_int_56_82 bl_int_55_82 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c83
+ bl_int_56_83 bl_int_55_83 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c84
+ bl_int_56_84 bl_int_55_84 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c85
+ bl_int_56_85 bl_int_55_85 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c86
+ bl_int_56_86 bl_int_55_86 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c87
+ bl_int_56_87 bl_int_55_87 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c88
+ bl_int_56_88 bl_int_55_88 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c89
+ bl_int_56_89 bl_int_55_89 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c90
+ bl_int_56_90 bl_int_55_90 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c91
+ bl_int_56_91 bl_int_55_91 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c92
+ bl_int_56_92 bl_int_55_92 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c93
+ bl_int_56_93 bl_int_55_93 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c94
+ bl_int_56_94 bl_int_55_94 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c95
+ bl_int_56_95 bl_int_55_95 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c96
+ bl_int_56_96 bl_int_55_96 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c97
+ bl_int_56_97 bl_int_55_97 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c98
+ bl_int_56_98 bl_int_55_98 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c99
+ bl_int_56_99 bl_int_55_99 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c100
+ bl_int_56_100 bl_int_55_100 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c101
+ bl_int_56_101 bl_int_55_101 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c102
+ bl_int_56_102 bl_int_55_102 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c103
+ bl_int_56_103 bl_int_55_103 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c104
+ bl_int_56_104 bl_int_55_104 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c105
+ bl_int_56_105 bl_int_55_105 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c106
+ bl_int_56_106 bl_int_55_106 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c107
+ bl_int_56_107 bl_int_55_107 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c108
+ bl_int_56_108 bl_int_55_108 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c109
+ bl_int_56_109 bl_int_55_109 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c110
+ bl_int_56_110 bl_int_55_110 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c111
+ bl_int_56_111 bl_int_55_111 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c112
+ bl_int_56_112 bl_int_55_112 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c113
+ bl_int_56_113 bl_int_55_113 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c114
+ bl_int_56_114 bl_int_55_114 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c115
+ bl_int_56_115 bl_int_55_115 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c116
+ bl_int_56_116 bl_int_55_116 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c117
+ bl_int_56_117 bl_int_55_117 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c118
+ bl_int_56_118 bl_int_55_118 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c119
+ bl_int_56_119 bl_int_55_119 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c120
+ bl_int_56_120 bl_int_55_120 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c121
+ bl_int_56_121 bl_int_55_121 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c122
+ bl_int_56_122 bl_int_55_122 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c123
+ bl_int_56_123 bl_int_55_123 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c124
+ bl_int_56_124 bl_int_55_124 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c125
+ bl_int_56_125 bl_int_55_125 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c126
+ bl_int_56_126 bl_int_55_126 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c127
+ bl_int_56_127 bl_int_55_127 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c128
+ bl_int_56_128 bl_int_55_128 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c129
+ bl_int_56_129 bl_int_55_129 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c130
+ bl_int_56_130 bl_int_55_130 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c131
+ bl_int_56_131 bl_int_55_131 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c132
+ bl_int_56_132 bl_int_55_132 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c133
+ bl_int_56_133 bl_int_55_133 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c134
+ bl_int_56_134 bl_int_55_134 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c135
+ bl_int_56_135 bl_int_55_135 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c136
+ bl_int_56_136 bl_int_55_136 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c137
+ bl_int_56_137 bl_int_55_137 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c138
+ bl_int_56_138 bl_int_55_138 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c139
+ bl_int_56_139 bl_int_55_139 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c140
+ bl_int_56_140 bl_int_55_140 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c141
+ bl_int_56_141 bl_int_55_141 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c142
+ bl_int_56_142 bl_int_55_142 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c143
+ bl_int_56_143 bl_int_55_143 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c144
+ bl_int_56_144 bl_int_55_144 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c145
+ bl_int_56_145 bl_int_55_145 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c146
+ bl_int_56_146 bl_int_55_146 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c147
+ bl_int_56_147 bl_int_55_147 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c148
+ bl_int_56_148 bl_int_55_148 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c149
+ bl_int_56_149 bl_int_55_149 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c150
+ bl_int_56_150 bl_int_55_150 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c151
+ bl_int_56_151 bl_int_55_151 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c152
+ bl_int_56_152 bl_int_55_152 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c153
+ bl_int_56_153 bl_int_55_153 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c154
+ bl_int_56_154 bl_int_55_154 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c155
+ bl_int_56_155 bl_int_55_155 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c156
+ bl_int_56_156 bl_int_55_156 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c157
+ bl_int_56_157 bl_int_55_157 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c158
+ bl_int_56_158 bl_int_55_158 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c159
+ bl_int_56_159 bl_int_55_159 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c160
+ bl_int_56_160 bl_int_55_160 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c161
+ bl_int_56_161 bl_int_55_161 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c162
+ bl_int_56_162 bl_int_55_162 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c163
+ bl_int_56_163 bl_int_55_163 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c164
+ bl_int_56_164 bl_int_55_164 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c165
+ bl_int_56_165 bl_int_55_165 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c166
+ bl_int_56_166 bl_int_55_166 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c167
+ bl_int_56_167 bl_int_55_167 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c168
+ bl_int_56_168 bl_int_55_168 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c169
+ bl_int_56_169 bl_int_55_169 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c170
+ bl_int_56_170 bl_int_55_170 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c171
+ bl_int_56_171 bl_int_55_171 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c172
+ bl_int_56_172 bl_int_55_172 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c173
+ bl_int_56_173 bl_int_55_173 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c174
+ bl_int_56_174 bl_int_55_174 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c175
+ bl_int_56_175 bl_int_55_175 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c176
+ bl_int_56_176 bl_int_55_176 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c177
+ bl_int_56_177 bl_int_55_177 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c178
+ bl_int_56_178 bl_int_55_178 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c179
+ bl_int_56_179 bl_int_55_179 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c180
+ bl_int_56_180 bl_int_55_180 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c181
+ bl_int_56_181 bl_int_55_181 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c182
+ bl_int_56_182 bl_int_55_182 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r56_c183
+ bl_int_56_183 bl_int_55_183 wl_0_56 gnd
+ sram_rom_base_one_cell
Xbit_r57_c0
+ bl_int_57_0 bl_int_56_0 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c1
+ bl_int_57_1 bl_int_56_1 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c2
+ bl_int_57_2 bl_int_56_2 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c3
+ bl_int_57_3 bl_int_56_3 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c4
+ bl_int_57_4 bl_int_56_4 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c5
+ bl_int_57_5 bl_int_56_5 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c6
+ bl_int_57_6 bl_int_56_6 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c7
+ bl_int_57_7 bl_int_56_7 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c8
+ bl_int_57_8 bl_int_56_8 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c9
+ bl_int_57_9 bl_int_56_9 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c10
+ bl_int_57_10 bl_int_56_10 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c11
+ bl_int_57_11 bl_int_56_11 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c12
+ bl_int_57_12 bl_int_56_12 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c13
+ bl_int_57_13 bl_int_56_13 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c14
+ bl_int_57_14 bl_int_56_14 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c15
+ bl_int_57_15 bl_int_56_15 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c16
+ bl_int_57_16 bl_int_56_16 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c17
+ bl_int_57_17 bl_int_56_17 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c18
+ bl_int_57_18 bl_int_56_18 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c19
+ bl_int_57_19 bl_int_56_19 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c20
+ bl_int_57_20 bl_int_56_20 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c21
+ bl_int_57_21 bl_int_56_21 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c22
+ bl_int_57_22 bl_int_56_22 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c23
+ bl_int_57_23 bl_int_56_23 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c24
+ bl_int_57_24 bl_int_56_24 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c25
+ bl_int_57_25 bl_int_56_25 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c26
+ bl_int_57_26 bl_int_56_26 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c27
+ bl_int_57_27 bl_int_56_27 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c28
+ bl_int_57_28 bl_int_56_28 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c29
+ bl_int_57_29 bl_int_56_29 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c30
+ bl_int_57_30 bl_int_56_30 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c31
+ bl_int_57_31 bl_int_56_31 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c32
+ bl_int_57_32 bl_int_56_32 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c33
+ bl_int_57_33 bl_int_56_33 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c34
+ bl_int_57_34 bl_int_56_34 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c35
+ bl_int_57_35 bl_int_56_35 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c36
+ bl_int_57_36 bl_int_56_36 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c37
+ bl_int_57_37 bl_int_56_37 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c38
+ bl_int_57_38 bl_int_56_38 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c39
+ bl_int_57_39 bl_int_56_39 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c40
+ bl_int_57_40 bl_int_56_40 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c41
+ bl_int_57_41 bl_int_56_41 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c42
+ bl_int_57_42 bl_int_56_42 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c43
+ bl_int_57_43 bl_int_56_43 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c44
+ bl_int_57_44 bl_int_56_44 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c45
+ bl_int_57_45 bl_int_56_45 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c46
+ bl_int_57_46 bl_int_56_46 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c47
+ bl_int_57_47 bl_int_56_47 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c48
+ bl_int_57_48 bl_int_56_48 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c49
+ bl_int_57_49 bl_int_56_49 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c50
+ bl_int_57_50 bl_int_56_50 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c51
+ bl_int_57_51 bl_int_56_51 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c52
+ bl_int_57_52 bl_int_56_52 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c53
+ bl_int_57_53 bl_int_56_53 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c54
+ bl_int_57_54 bl_int_56_54 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c55
+ bl_int_57_55 bl_int_56_55 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c56
+ bl_int_57_56 bl_int_56_56 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c57
+ bl_int_57_57 bl_int_56_57 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c58
+ bl_int_57_58 bl_int_56_58 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c59
+ bl_int_57_59 bl_int_56_59 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c60
+ bl_int_57_60 bl_int_56_60 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c61
+ bl_int_57_61 bl_int_56_61 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c62
+ bl_int_57_62 bl_int_56_62 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c63
+ bl_int_57_63 bl_int_56_63 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c64
+ bl_int_57_64 bl_int_56_64 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c65
+ bl_int_57_65 bl_int_56_65 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c66
+ bl_int_57_66 bl_int_56_66 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c67
+ bl_int_57_67 bl_int_56_67 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c68
+ bl_int_57_68 bl_int_56_68 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c69
+ bl_int_57_69 bl_int_56_69 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c70
+ bl_int_57_70 bl_int_56_70 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c71
+ bl_int_57_71 bl_int_56_71 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c72
+ bl_int_57_72 bl_int_56_72 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c73
+ bl_int_57_73 bl_int_56_73 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c74
+ bl_int_57_74 bl_int_56_74 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c75
+ bl_int_57_75 bl_int_56_75 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c76
+ bl_int_57_76 bl_int_56_76 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c77
+ bl_int_57_77 bl_int_56_77 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c78
+ bl_int_57_78 bl_int_56_78 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c79
+ bl_int_57_79 bl_int_56_79 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c80
+ bl_int_57_80 bl_int_56_80 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c81
+ bl_int_57_81 bl_int_56_81 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c82
+ bl_int_57_82 bl_int_56_82 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c83
+ bl_int_57_83 bl_int_56_83 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c84
+ bl_int_57_84 bl_int_56_84 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c85
+ bl_int_57_85 bl_int_56_85 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c86
+ bl_int_57_86 bl_int_56_86 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c87
+ bl_int_57_87 bl_int_56_87 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c88
+ bl_int_57_88 bl_int_56_88 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c89
+ bl_int_57_89 bl_int_56_89 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c90
+ bl_int_57_90 bl_int_56_90 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c91
+ bl_int_57_91 bl_int_56_91 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c92
+ bl_int_57_92 bl_int_56_92 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c93
+ bl_int_57_93 bl_int_56_93 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c94
+ bl_int_57_94 bl_int_56_94 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c95
+ bl_int_57_95 bl_int_56_95 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c96
+ bl_int_57_96 bl_int_56_96 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c97
+ bl_int_57_97 bl_int_56_97 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c98
+ bl_int_57_98 bl_int_56_98 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c99
+ bl_int_57_99 bl_int_56_99 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c100
+ bl_int_57_100 bl_int_56_100 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c101
+ bl_int_57_101 bl_int_56_101 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c102
+ bl_int_57_102 bl_int_56_102 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c103
+ bl_int_57_103 bl_int_56_103 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c104
+ bl_int_57_104 bl_int_56_104 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c105
+ bl_int_57_105 bl_int_56_105 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c106
+ bl_int_57_106 bl_int_56_106 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c107
+ bl_int_57_107 bl_int_56_107 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c108
+ bl_int_57_108 bl_int_56_108 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c109
+ bl_int_57_109 bl_int_56_109 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c110
+ bl_int_57_110 bl_int_56_110 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c111
+ bl_int_57_111 bl_int_56_111 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c112
+ bl_int_57_112 bl_int_56_112 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c113
+ bl_int_57_113 bl_int_56_113 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c114
+ bl_int_57_114 bl_int_56_114 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c115
+ bl_int_57_115 bl_int_56_115 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c116
+ bl_int_57_116 bl_int_56_116 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c117
+ bl_int_57_117 bl_int_56_117 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c118
+ bl_int_57_118 bl_int_56_118 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c119
+ bl_int_57_119 bl_int_56_119 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c120
+ bl_int_57_120 bl_int_56_120 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c121
+ bl_int_57_121 bl_int_56_121 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c122
+ bl_int_57_122 bl_int_56_122 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c123
+ bl_int_57_123 bl_int_56_123 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c124
+ bl_int_57_124 bl_int_56_124 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c125
+ bl_int_57_125 bl_int_56_125 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c126
+ bl_int_57_126 bl_int_56_126 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c127
+ bl_int_57_127 bl_int_56_127 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c128
+ bl_int_57_128 bl_int_56_128 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c129
+ bl_int_57_129 bl_int_56_129 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c130
+ bl_int_57_130 bl_int_56_130 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c131
+ bl_int_57_131 bl_int_56_131 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c132
+ bl_int_57_132 bl_int_56_132 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c133
+ bl_int_57_133 bl_int_56_133 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c134
+ bl_int_57_134 bl_int_56_134 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c135
+ bl_int_57_135 bl_int_56_135 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c136
+ bl_int_57_136 bl_int_56_136 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c137
+ bl_int_57_137 bl_int_56_137 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c138
+ bl_int_57_138 bl_int_56_138 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c139
+ bl_int_57_139 bl_int_56_139 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c140
+ bl_int_57_140 bl_int_56_140 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c141
+ bl_int_57_141 bl_int_56_141 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c142
+ bl_int_57_142 bl_int_56_142 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c143
+ bl_int_57_143 bl_int_56_143 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c144
+ bl_int_57_144 bl_int_56_144 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c145
+ bl_int_57_145 bl_int_56_145 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c146
+ bl_int_57_146 bl_int_56_146 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c147
+ bl_int_57_147 bl_int_56_147 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c148
+ bl_int_57_148 bl_int_56_148 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c149
+ bl_int_57_149 bl_int_56_149 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c150
+ bl_int_57_150 bl_int_56_150 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c151
+ bl_int_57_151 bl_int_56_151 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c152
+ bl_int_57_152 bl_int_56_152 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c153
+ bl_int_57_153 bl_int_56_153 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c154
+ bl_int_57_154 bl_int_56_154 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c155
+ bl_int_57_155 bl_int_56_155 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c156
+ bl_int_57_156 bl_int_56_156 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c157
+ bl_int_57_157 bl_int_56_157 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c158
+ bl_int_57_158 bl_int_56_158 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c159
+ bl_int_57_159 bl_int_56_159 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c160
+ bl_int_57_160 bl_int_56_160 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c161
+ bl_int_57_161 bl_int_56_161 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c162
+ bl_int_57_162 bl_int_56_162 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c163
+ bl_int_57_163 bl_int_56_163 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c164
+ bl_int_57_164 bl_int_56_164 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c165
+ bl_int_57_165 bl_int_56_165 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c166
+ bl_int_57_166 bl_int_56_166 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c167
+ bl_int_57_167 bl_int_56_167 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c168
+ bl_int_57_168 bl_int_56_168 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c169
+ bl_int_57_169 bl_int_56_169 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c170
+ bl_int_57_170 bl_int_56_170 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c171
+ bl_int_57_171 bl_int_56_171 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c172
+ bl_int_57_172 bl_int_56_172 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c173
+ bl_int_57_173 bl_int_56_173 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c174
+ bl_int_57_174 bl_int_56_174 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c175
+ bl_int_57_175 bl_int_56_175 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c176
+ bl_int_57_176 bl_int_56_176 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c177
+ bl_int_57_177 bl_int_56_177 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c178
+ bl_int_57_178 bl_int_56_178 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c179
+ bl_int_57_179 bl_int_56_179 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c180
+ bl_int_57_180 bl_int_56_180 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c181
+ bl_int_57_181 bl_int_56_181 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c182
+ bl_int_57_182 bl_int_56_182 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r57_c183
+ bl_int_57_183 bl_int_56_183 wl_0_57 gnd
+ sram_rom_base_one_cell
Xbit_r58_c0
+ bl_int_58_0 bl_int_57_0 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c1
+ bl_int_58_1 bl_int_57_1 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c2
+ bl_int_58_2 bl_int_57_2 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c3
+ bl_int_58_3 bl_int_57_3 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c4
+ bl_int_58_4 bl_int_57_4 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c5
+ bl_int_58_5 bl_int_57_5 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c6
+ bl_int_58_6 bl_int_57_6 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c7
+ bl_int_58_7 bl_int_57_7 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c8
+ bl_int_58_8 bl_int_57_8 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c9
+ bl_int_58_9 bl_int_57_9 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c10
+ bl_int_58_10 bl_int_57_10 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c11
+ bl_int_58_11 bl_int_57_11 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c12
+ bl_int_58_12 bl_int_57_12 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c13
+ bl_int_58_13 bl_int_57_13 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c14
+ bl_int_58_14 bl_int_57_14 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c15
+ bl_int_58_15 bl_int_57_15 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c16
+ bl_int_58_16 bl_int_57_16 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c17
+ bl_int_58_17 bl_int_57_17 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c18
+ bl_int_58_18 bl_int_57_18 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c19
+ bl_int_58_19 bl_int_57_19 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c20
+ bl_int_58_20 bl_int_57_20 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c21
+ bl_int_58_21 bl_int_57_21 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c22
+ bl_int_58_22 bl_int_57_22 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c23
+ bl_int_58_23 bl_int_57_23 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c24
+ bl_int_58_24 bl_int_57_24 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c25
+ bl_int_58_25 bl_int_57_25 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c26
+ bl_int_58_26 bl_int_57_26 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c27
+ bl_int_58_27 bl_int_57_27 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c28
+ bl_int_58_28 bl_int_57_28 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c29
+ bl_int_58_29 bl_int_57_29 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c30
+ bl_int_58_30 bl_int_57_30 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c31
+ bl_int_58_31 bl_int_57_31 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c32
+ bl_int_58_32 bl_int_57_32 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c33
+ bl_int_58_33 bl_int_57_33 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c34
+ bl_int_58_34 bl_int_57_34 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c35
+ bl_int_58_35 bl_int_57_35 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c36
+ bl_int_58_36 bl_int_57_36 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c37
+ bl_int_58_37 bl_int_57_37 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c38
+ bl_int_58_38 bl_int_57_38 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c39
+ bl_int_58_39 bl_int_57_39 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c40
+ bl_int_58_40 bl_int_57_40 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c41
+ bl_int_58_41 bl_int_57_41 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c42
+ bl_int_58_42 bl_int_57_42 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c43
+ bl_int_58_43 bl_int_57_43 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c44
+ bl_int_58_44 bl_int_57_44 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c45
+ bl_int_58_45 bl_int_57_45 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c46
+ bl_int_58_46 bl_int_57_46 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c47
+ bl_int_58_47 bl_int_57_47 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c48
+ bl_int_58_48 bl_int_57_48 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c49
+ bl_int_58_49 bl_int_57_49 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c50
+ bl_int_58_50 bl_int_57_50 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c51
+ bl_int_58_51 bl_int_57_51 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c52
+ bl_int_58_52 bl_int_57_52 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c53
+ bl_int_58_53 bl_int_57_53 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c54
+ bl_int_58_54 bl_int_57_54 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c55
+ bl_int_58_55 bl_int_57_55 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c56
+ bl_int_58_56 bl_int_57_56 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c57
+ bl_int_58_57 bl_int_57_57 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c58
+ bl_int_58_58 bl_int_57_58 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c59
+ bl_int_58_59 bl_int_57_59 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c60
+ bl_int_58_60 bl_int_57_60 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c61
+ bl_int_58_61 bl_int_57_61 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c62
+ bl_int_58_62 bl_int_57_62 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c63
+ bl_int_58_63 bl_int_57_63 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c64
+ bl_int_58_64 bl_int_57_64 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c65
+ bl_int_58_65 bl_int_57_65 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c66
+ bl_int_58_66 bl_int_57_66 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c67
+ bl_int_58_67 bl_int_57_67 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c68
+ bl_int_58_68 bl_int_57_68 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c69
+ bl_int_58_69 bl_int_57_69 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c70
+ bl_int_58_70 bl_int_57_70 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c71
+ bl_int_58_71 bl_int_57_71 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c72
+ bl_int_58_72 bl_int_57_72 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c73
+ bl_int_58_73 bl_int_57_73 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c74
+ bl_int_58_74 bl_int_57_74 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c75
+ bl_int_58_75 bl_int_57_75 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c76
+ bl_int_58_76 bl_int_57_76 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c77
+ bl_int_58_77 bl_int_57_77 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c78
+ bl_int_58_78 bl_int_57_78 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c79
+ bl_int_58_79 bl_int_57_79 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c80
+ bl_int_58_80 bl_int_57_80 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c81
+ bl_int_58_81 bl_int_57_81 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c82
+ bl_int_58_82 bl_int_57_82 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c83
+ bl_int_58_83 bl_int_57_83 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c84
+ bl_int_58_84 bl_int_57_84 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c85
+ bl_int_58_85 bl_int_57_85 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c86
+ bl_int_58_86 bl_int_57_86 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c87
+ bl_int_58_87 bl_int_57_87 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c88
+ bl_int_58_88 bl_int_57_88 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c89
+ bl_int_58_89 bl_int_57_89 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c90
+ bl_int_58_90 bl_int_57_90 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c91
+ bl_int_58_91 bl_int_57_91 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c92
+ bl_int_58_92 bl_int_57_92 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c93
+ bl_int_58_93 bl_int_57_93 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c94
+ bl_int_58_94 bl_int_57_94 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c95
+ bl_int_58_95 bl_int_57_95 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c96
+ bl_int_58_96 bl_int_57_96 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c97
+ bl_int_58_97 bl_int_57_97 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c98
+ bl_int_58_98 bl_int_57_98 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c99
+ bl_int_58_99 bl_int_57_99 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c100
+ bl_int_58_100 bl_int_57_100 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c101
+ bl_int_58_101 bl_int_57_101 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c102
+ bl_int_58_102 bl_int_57_102 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c103
+ bl_int_58_103 bl_int_57_103 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c104
+ bl_int_58_104 bl_int_57_104 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c105
+ bl_int_58_105 bl_int_57_105 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c106
+ bl_int_58_106 bl_int_57_106 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c107
+ bl_int_58_107 bl_int_57_107 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c108
+ bl_int_58_108 bl_int_57_108 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c109
+ bl_int_58_109 bl_int_57_109 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c110
+ bl_int_58_110 bl_int_57_110 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c111
+ bl_int_58_111 bl_int_57_111 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c112
+ bl_int_58_112 bl_int_57_112 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c113
+ bl_int_58_113 bl_int_57_113 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c114
+ bl_int_58_114 bl_int_57_114 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c115
+ bl_int_58_115 bl_int_57_115 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c116
+ bl_int_58_116 bl_int_57_116 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c117
+ bl_int_58_117 bl_int_57_117 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c118
+ bl_int_58_118 bl_int_57_118 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c119
+ bl_int_58_119 bl_int_57_119 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c120
+ bl_int_58_120 bl_int_57_120 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c121
+ bl_int_58_121 bl_int_57_121 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c122
+ bl_int_58_122 bl_int_57_122 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c123
+ bl_int_58_123 bl_int_57_123 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c124
+ bl_int_58_124 bl_int_57_124 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c125
+ bl_int_58_125 bl_int_57_125 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c126
+ bl_int_58_126 bl_int_57_126 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c127
+ bl_int_58_127 bl_int_57_127 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c128
+ bl_int_58_128 bl_int_57_128 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c129
+ bl_int_58_129 bl_int_57_129 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c130
+ bl_int_58_130 bl_int_57_130 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c131
+ bl_int_58_131 bl_int_57_131 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c132
+ bl_int_58_132 bl_int_57_132 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c133
+ bl_int_58_133 bl_int_57_133 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c134
+ bl_int_58_134 bl_int_57_134 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c135
+ bl_int_58_135 bl_int_57_135 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c136
+ bl_int_58_136 bl_int_57_136 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c137
+ bl_int_58_137 bl_int_57_137 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c138
+ bl_int_58_138 bl_int_57_138 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c139
+ bl_int_58_139 bl_int_57_139 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c140
+ bl_int_58_140 bl_int_57_140 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c141
+ bl_int_58_141 bl_int_57_141 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c142
+ bl_int_58_142 bl_int_57_142 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c143
+ bl_int_58_143 bl_int_57_143 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c144
+ bl_int_58_144 bl_int_57_144 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c145
+ bl_int_58_145 bl_int_57_145 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c146
+ bl_int_58_146 bl_int_57_146 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c147
+ bl_int_58_147 bl_int_57_147 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c148
+ bl_int_58_148 bl_int_57_148 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c149
+ bl_int_58_149 bl_int_57_149 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c150
+ bl_int_58_150 bl_int_57_150 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c151
+ bl_int_58_151 bl_int_57_151 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c152
+ bl_int_58_152 bl_int_57_152 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c153
+ bl_int_58_153 bl_int_57_153 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c154
+ bl_int_58_154 bl_int_57_154 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c155
+ bl_int_58_155 bl_int_57_155 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c156
+ bl_int_58_156 bl_int_57_156 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c157
+ bl_int_58_157 bl_int_57_157 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c158
+ bl_int_58_158 bl_int_57_158 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c159
+ bl_int_58_159 bl_int_57_159 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c160
+ bl_int_58_160 bl_int_57_160 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c161
+ bl_int_58_161 bl_int_57_161 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c162
+ bl_int_58_162 bl_int_57_162 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c163
+ bl_int_58_163 bl_int_57_163 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c164
+ bl_int_58_164 bl_int_57_164 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c165
+ bl_int_58_165 bl_int_57_165 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c166
+ bl_int_58_166 bl_int_57_166 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c167
+ bl_int_58_167 bl_int_57_167 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c168
+ bl_int_58_168 bl_int_57_168 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c169
+ bl_int_58_169 bl_int_57_169 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c170
+ bl_int_58_170 bl_int_57_170 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c171
+ bl_int_58_171 bl_int_57_171 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c172
+ bl_int_58_172 bl_int_57_172 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c173
+ bl_int_58_173 bl_int_57_173 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c174
+ bl_int_58_174 bl_int_57_174 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c175
+ bl_int_58_175 bl_int_57_175 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c176
+ bl_int_58_176 bl_int_57_176 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c177
+ bl_int_58_177 bl_int_57_177 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c178
+ bl_int_58_178 bl_int_57_178 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c179
+ bl_int_58_179 bl_int_57_179 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c180
+ bl_int_58_180 bl_int_57_180 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c181
+ bl_int_58_181 bl_int_57_181 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c182
+ bl_int_58_182 bl_int_57_182 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r58_c183
+ bl_int_58_183 bl_int_57_183 wl_0_58 gnd
+ sram_rom_base_one_cell
Xbit_r59_c0
+ bl_int_59_0 bl_int_58_0 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c1
+ bl_int_59_1 bl_int_58_1 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c2
+ bl_int_59_2 bl_int_58_2 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c3
+ bl_int_59_3 bl_int_58_3 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c4
+ bl_int_59_4 bl_int_58_4 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c5
+ bl_int_59_5 bl_int_58_5 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c6
+ bl_int_59_6 bl_int_58_6 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c7
+ bl_int_59_7 bl_int_58_7 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c8
+ bl_int_59_8 bl_int_58_8 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c9
+ bl_int_59_9 bl_int_58_9 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c10
+ bl_int_59_10 bl_int_58_10 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c11
+ bl_int_59_11 bl_int_58_11 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c12
+ bl_int_59_12 bl_int_58_12 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c13
+ bl_int_59_13 bl_int_58_13 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c14
+ bl_int_59_14 bl_int_58_14 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c15
+ bl_int_59_15 bl_int_58_15 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c16
+ bl_int_59_16 bl_int_58_16 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c17
+ bl_int_59_17 bl_int_58_17 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c18
+ bl_int_59_18 bl_int_58_18 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c19
+ bl_int_59_19 bl_int_58_19 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c20
+ bl_int_59_20 bl_int_58_20 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c21
+ bl_int_59_21 bl_int_58_21 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c22
+ bl_int_59_22 bl_int_58_22 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c23
+ bl_int_59_23 bl_int_58_23 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c24
+ bl_int_59_24 bl_int_58_24 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c25
+ bl_int_59_25 bl_int_58_25 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c26
+ bl_int_59_26 bl_int_58_26 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c27
+ bl_int_59_27 bl_int_58_27 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c28
+ bl_int_59_28 bl_int_58_28 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c29
+ bl_int_59_29 bl_int_58_29 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c30
+ bl_int_59_30 bl_int_58_30 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c31
+ bl_int_59_31 bl_int_58_31 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c32
+ bl_int_59_32 bl_int_58_32 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c33
+ bl_int_59_33 bl_int_58_33 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c34
+ bl_int_59_34 bl_int_58_34 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c35
+ bl_int_59_35 bl_int_58_35 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c36
+ bl_int_59_36 bl_int_58_36 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c37
+ bl_int_59_37 bl_int_58_37 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c38
+ bl_int_59_38 bl_int_58_38 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c39
+ bl_int_59_39 bl_int_58_39 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c40
+ bl_int_59_40 bl_int_58_40 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c41
+ bl_int_59_41 bl_int_58_41 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c42
+ bl_int_59_42 bl_int_58_42 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c43
+ bl_int_59_43 bl_int_58_43 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c44
+ bl_int_59_44 bl_int_58_44 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c45
+ bl_int_59_45 bl_int_58_45 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c46
+ bl_int_59_46 bl_int_58_46 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c47
+ bl_int_59_47 bl_int_58_47 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c48
+ bl_int_59_48 bl_int_58_48 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c49
+ bl_int_59_49 bl_int_58_49 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c50
+ bl_int_59_50 bl_int_58_50 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c51
+ bl_int_59_51 bl_int_58_51 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c52
+ bl_int_59_52 bl_int_58_52 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c53
+ bl_int_59_53 bl_int_58_53 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c54
+ bl_int_59_54 bl_int_58_54 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c55
+ bl_int_59_55 bl_int_58_55 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c56
+ bl_int_59_56 bl_int_58_56 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c57
+ bl_int_59_57 bl_int_58_57 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c58
+ bl_int_59_58 bl_int_58_58 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c59
+ bl_int_59_59 bl_int_58_59 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c60
+ bl_int_59_60 bl_int_58_60 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c61
+ bl_int_59_61 bl_int_58_61 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c62
+ bl_int_59_62 bl_int_58_62 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c63
+ bl_int_59_63 bl_int_58_63 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c64
+ bl_int_59_64 bl_int_58_64 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c65
+ bl_int_59_65 bl_int_58_65 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c66
+ bl_int_59_66 bl_int_58_66 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c67
+ bl_int_59_67 bl_int_58_67 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c68
+ bl_int_59_68 bl_int_58_68 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c69
+ bl_int_59_69 bl_int_58_69 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c70
+ bl_int_59_70 bl_int_58_70 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c71
+ bl_int_59_71 bl_int_58_71 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c72
+ bl_int_59_72 bl_int_58_72 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c73
+ bl_int_59_73 bl_int_58_73 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c74
+ bl_int_59_74 bl_int_58_74 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c75
+ bl_int_59_75 bl_int_58_75 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c76
+ bl_int_59_76 bl_int_58_76 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c77
+ bl_int_59_77 bl_int_58_77 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c78
+ bl_int_59_78 bl_int_58_78 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c79
+ bl_int_59_79 bl_int_58_79 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c80
+ bl_int_59_80 bl_int_58_80 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c81
+ bl_int_59_81 bl_int_58_81 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c82
+ bl_int_59_82 bl_int_58_82 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c83
+ bl_int_59_83 bl_int_58_83 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c84
+ bl_int_59_84 bl_int_58_84 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c85
+ bl_int_59_85 bl_int_58_85 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c86
+ bl_int_59_86 bl_int_58_86 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c87
+ bl_int_59_87 bl_int_58_87 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c88
+ bl_int_59_88 bl_int_58_88 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c89
+ bl_int_59_89 bl_int_58_89 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c90
+ bl_int_59_90 bl_int_58_90 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c91
+ bl_int_59_91 bl_int_58_91 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c92
+ bl_int_59_92 bl_int_58_92 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c93
+ bl_int_59_93 bl_int_58_93 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c94
+ bl_int_59_94 bl_int_58_94 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c95
+ bl_int_59_95 bl_int_58_95 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c96
+ bl_int_59_96 bl_int_58_96 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c97
+ bl_int_59_97 bl_int_58_97 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c98
+ bl_int_59_98 bl_int_58_98 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c99
+ bl_int_59_99 bl_int_58_99 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c100
+ bl_int_59_100 bl_int_58_100 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c101
+ bl_int_59_101 bl_int_58_101 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c102
+ bl_int_59_102 bl_int_58_102 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c103
+ bl_int_59_103 bl_int_58_103 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c104
+ bl_int_59_104 bl_int_58_104 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c105
+ bl_int_59_105 bl_int_58_105 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c106
+ bl_int_59_106 bl_int_58_106 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c107
+ bl_int_59_107 bl_int_58_107 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c108
+ bl_int_59_108 bl_int_58_108 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c109
+ bl_int_59_109 bl_int_58_109 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c110
+ bl_int_59_110 bl_int_58_110 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c111
+ bl_int_59_111 bl_int_58_111 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c112
+ bl_int_59_112 bl_int_58_112 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c113
+ bl_int_59_113 bl_int_58_113 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c114
+ bl_int_59_114 bl_int_58_114 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c115
+ bl_int_59_115 bl_int_58_115 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c116
+ bl_int_59_116 bl_int_58_116 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c117
+ bl_int_59_117 bl_int_58_117 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c118
+ bl_int_59_118 bl_int_58_118 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c119
+ bl_int_59_119 bl_int_58_119 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c120
+ bl_int_59_120 bl_int_58_120 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c121
+ bl_int_59_121 bl_int_58_121 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c122
+ bl_int_59_122 bl_int_58_122 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c123
+ bl_int_59_123 bl_int_58_123 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c124
+ bl_int_59_124 bl_int_58_124 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c125
+ bl_int_59_125 bl_int_58_125 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c126
+ bl_int_59_126 bl_int_58_126 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c127
+ bl_int_59_127 bl_int_58_127 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c128
+ bl_int_59_128 bl_int_58_128 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c129
+ bl_int_59_129 bl_int_58_129 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c130
+ bl_int_59_130 bl_int_58_130 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c131
+ bl_int_59_131 bl_int_58_131 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c132
+ bl_int_59_132 bl_int_58_132 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c133
+ bl_int_59_133 bl_int_58_133 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c134
+ bl_int_59_134 bl_int_58_134 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c135
+ bl_int_59_135 bl_int_58_135 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c136
+ bl_int_59_136 bl_int_58_136 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c137
+ bl_int_59_137 bl_int_58_137 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c138
+ bl_int_59_138 bl_int_58_138 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c139
+ bl_int_59_139 bl_int_58_139 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c140
+ bl_int_59_140 bl_int_58_140 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c141
+ bl_int_59_141 bl_int_58_141 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c142
+ bl_int_59_142 bl_int_58_142 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c143
+ bl_int_59_143 bl_int_58_143 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c144
+ bl_int_59_144 bl_int_58_144 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c145
+ bl_int_59_145 bl_int_58_145 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c146
+ bl_int_59_146 bl_int_58_146 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c147
+ bl_int_59_147 bl_int_58_147 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c148
+ bl_int_59_148 bl_int_58_148 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c149
+ bl_int_59_149 bl_int_58_149 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c150
+ bl_int_59_150 bl_int_58_150 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c151
+ bl_int_59_151 bl_int_58_151 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c152
+ bl_int_59_152 bl_int_58_152 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c153
+ bl_int_59_153 bl_int_58_153 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c154
+ bl_int_59_154 bl_int_58_154 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c155
+ bl_int_59_155 bl_int_58_155 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c156
+ bl_int_59_156 bl_int_58_156 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c157
+ bl_int_59_157 bl_int_58_157 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c158
+ bl_int_59_158 bl_int_58_158 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c159
+ bl_int_59_159 bl_int_58_159 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c160
+ bl_int_59_160 bl_int_58_160 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c161
+ bl_int_59_161 bl_int_58_161 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c162
+ bl_int_59_162 bl_int_58_162 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c163
+ bl_int_59_163 bl_int_58_163 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c164
+ bl_int_59_164 bl_int_58_164 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c165
+ bl_int_59_165 bl_int_58_165 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c166
+ bl_int_59_166 bl_int_58_166 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c167
+ bl_int_59_167 bl_int_58_167 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c168
+ bl_int_59_168 bl_int_58_168 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c169
+ bl_int_59_169 bl_int_58_169 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c170
+ bl_int_59_170 bl_int_58_170 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c171
+ bl_int_59_171 bl_int_58_171 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c172
+ bl_int_59_172 bl_int_58_172 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c173
+ bl_int_59_173 bl_int_58_173 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c174
+ bl_int_59_174 bl_int_58_174 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c175
+ bl_int_59_175 bl_int_58_175 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c176
+ bl_int_59_176 bl_int_58_176 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c177
+ bl_int_59_177 bl_int_58_177 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c178
+ bl_int_59_178 bl_int_58_178 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c179
+ bl_int_59_179 bl_int_58_179 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c180
+ bl_int_59_180 bl_int_58_180 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c181
+ bl_int_59_181 bl_int_58_181 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c182
+ bl_int_59_182 bl_int_58_182 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r59_c183
+ bl_int_59_183 bl_int_58_183 wl_0_59 gnd
+ sram_rom_base_one_cell
Xbit_r60_c0
+ bl_int_60_0 bl_int_59_0 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c1
+ bl_int_60_1 bl_int_59_1 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c2
+ bl_int_60_2 bl_int_59_2 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c3
+ bl_int_60_3 bl_int_59_3 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c4
+ bl_int_60_4 bl_int_59_4 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c5
+ bl_int_60_5 bl_int_59_5 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c6
+ bl_int_60_6 bl_int_59_6 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c7
+ bl_int_60_7 bl_int_59_7 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c8
+ bl_int_60_8 bl_int_59_8 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c9
+ bl_int_60_9 bl_int_59_9 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c10
+ bl_int_60_10 bl_int_59_10 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c11
+ bl_int_60_11 bl_int_59_11 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c12
+ bl_int_60_12 bl_int_59_12 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c13
+ bl_int_60_13 bl_int_59_13 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c14
+ bl_int_60_14 bl_int_59_14 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c15
+ bl_int_60_15 bl_int_59_15 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c16
+ bl_int_60_16 bl_int_59_16 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c17
+ bl_int_60_17 bl_int_59_17 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c18
+ bl_int_60_18 bl_int_59_18 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c19
+ bl_int_60_19 bl_int_59_19 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c20
+ bl_int_60_20 bl_int_59_20 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c21
+ bl_int_60_21 bl_int_59_21 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c22
+ bl_int_60_22 bl_int_59_22 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c23
+ bl_int_60_23 bl_int_59_23 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c24
+ bl_int_60_24 bl_int_59_24 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c25
+ bl_int_60_25 bl_int_59_25 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c26
+ bl_int_60_26 bl_int_59_26 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c27
+ bl_int_60_27 bl_int_59_27 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c28
+ bl_int_60_28 bl_int_59_28 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c29
+ bl_int_60_29 bl_int_59_29 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c30
+ bl_int_60_30 bl_int_59_30 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c31
+ bl_int_60_31 bl_int_59_31 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c32
+ bl_int_60_32 bl_int_59_32 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c33
+ bl_int_60_33 bl_int_59_33 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c34
+ bl_int_60_34 bl_int_59_34 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c35
+ bl_int_60_35 bl_int_59_35 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c36
+ bl_int_60_36 bl_int_59_36 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c37
+ bl_int_60_37 bl_int_59_37 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c38
+ bl_int_60_38 bl_int_59_38 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c39
+ bl_int_60_39 bl_int_59_39 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c40
+ bl_int_60_40 bl_int_59_40 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c41
+ bl_int_60_41 bl_int_59_41 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c42
+ bl_int_60_42 bl_int_59_42 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c43
+ bl_int_60_43 bl_int_59_43 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c44
+ bl_int_60_44 bl_int_59_44 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c45
+ bl_int_60_45 bl_int_59_45 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c46
+ bl_int_60_46 bl_int_59_46 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c47
+ bl_int_60_47 bl_int_59_47 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c48
+ bl_int_60_48 bl_int_59_48 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c49
+ bl_int_60_49 bl_int_59_49 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c50
+ bl_int_60_50 bl_int_59_50 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c51
+ bl_int_60_51 bl_int_59_51 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c52
+ bl_int_60_52 bl_int_59_52 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c53
+ bl_int_60_53 bl_int_59_53 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c54
+ bl_int_60_54 bl_int_59_54 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c55
+ bl_int_60_55 bl_int_59_55 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c56
+ bl_int_60_56 bl_int_59_56 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c57
+ bl_int_60_57 bl_int_59_57 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c58
+ bl_int_60_58 bl_int_59_58 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c59
+ bl_int_60_59 bl_int_59_59 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c60
+ bl_int_60_60 bl_int_59_60 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c61
+ bl_int_60_61 bl_int_59_61 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c62
+ bl_int_60_62 bl_int_59_62 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c63
+ bl_int_60_63 bl_int_59_63 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c64
+ bl_int_60_64 bl_int_59_64 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c65
+ bl_int_60_65 bl_int_59_65 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c66
+ bl_int_60_66 bl_int_59_66 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c67
+ bl_int_60_67 bl_int_59_67 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c68
+ bl_int_60_68 bl_int_59_68 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c69
+ bl_int_60_69 bl_int_59_69 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c70
+ bl_int_60_70 bl_int_59_70 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c71
+ bl_int_60_71 bl_int_59_71 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c72
+ bl_int_60_72 bl_int_59_72 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c73
+ bl_int_60_73 bl_int_59_73 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c74
+ bl_int_60_74 bl_int_59_74 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c75
+ bl_int_60_75 bl_int_59_75 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c76
+ bl_int_60_76 bl_int_59_76 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c77
+ bl_int_60_77 bl_int_59_77 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c78
+ bl_int_60_78 bl_int_59_78 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c79
+ bl_int_60_79 bl_int_59_79 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c80
+ bl_int_60_80 bl_int_59_80 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c81
+ bl_int_60_81 bl_int_59_81 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c82
+ bl_int_60_82 bl_int_59_82 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c83
+ bl_int_60_83 bl_int_59_83 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c84
+ bl_int_60_84 bl_int_59_84 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c85
+ bl_int_60_85 bl_int_59_85 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c86
+ bl_int_60_86 bl_int_59_86 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c87
+ bl_int_60_87 bl_int_59_87 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c88
+ bl_int_60_88 bl_int_59_88 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c89
+ bl_int_60_89 bl_int_59_89 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c90
+ bl_int_60_90 bl_int_59_90 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c91
+ bl_int_60_91 bl_int_59_91 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c92
+ bl_int_60_92 bl_int_59_92 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c93
+ bl_int_60_93 bl_int_59_93 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c94
+ bl_int_60_94 bl_int_59_94 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c95
+ bl_int_60_95 bl_int_59_95 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c96
+ bl_int_60_96 bl_int_59_96 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c97
+ bl_int_60_97 bl_int_59_97 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c98
+ bl_int_60_98 bl_int_59_98 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c99
+ bl_int_60_99 bl_int_59_99 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c100
+ bl_int_60_100 bl_int_59_100 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c101
+ bl_int_60_101 bl_int_59_101 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c102
+ bl_int_60_102 bl_int_59_102 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c103
+ bl_int_60_103 bl_int_59_103 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c104
+ bl_int_60_104 bl_int_59_104 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c105
+ bl_int_60_105 bl_int_59_105 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c106
+ bl_int_60_106 bl_int_59_106 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c107
+ bl_int_60_107 bl_int_59_107 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c108
+ bl_int_60_108 bl_int_59_108 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c109
+ bl_int_60_109 bl_int_59_109 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c110
+ bl_int_60_110 bl_int_59_110 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c111
+ bl_int_60_111 bl_int_59_111 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c112
+ bl_int_60_112 bl_int_59_112 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c113
+ bl_int_60_113 bl_int_59_113 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c114
+ bl_int_60_114 bl_int_59_114 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c115
+ bl_int_60_115 bl_int_59_115 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c116
+ bl_int_60_116 bl_int_59_116 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c117
+ bl_int_60_117 bl_int_59_117 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c118
+ bl_int_60_118 bl_int_59_118 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c119
+ bl_int_60_119 bl_int_59_119 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c120
+ bl_int_60_120 bl_int_59_120 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c121
+ bl_int_60_121 bl_int_59_121 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c122
+ bl_int_60_122 bl_int_59_122 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c123
+ bl_int_60_123 bl_int_59_123 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c124
+ bl_int_60_124 bl_int_59_124 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c125
+ bl_int_60_125 bl_int_59_125 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c126
+ bl_int_60_126 bl_int_59_126 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c127
+ bl_int_60_127 bl_int_59_127 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c128
+ bl_int_60_128 bl_int_59_128 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c129
+ bl_int_60_129 bl_int_59_129 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c130
+ bl_int_60_130 bl_int_59_130 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c131
+ bl_int_60_131 bl_int_59_131 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c132
+ bl_int_60_132 bl_int_59_132 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c133
+ bl_int_60_133 bl_int_59_133 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c134
+ bl_int_60_134 bl_int_59_134 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c135
+ bl_int_60_135 bl_int_59_135 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c136
+ bl_int_60_136 bl_int_59_136 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c137
+ bl_int_60_137 bl_int_59_137 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c138
+ bl_int_60_138 bl_int_59_138 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c139
+ bl_int_60_139 bl_int_59_139 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c140
+ bl_int_60_140 bl_int_59_140 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c141
+ bl_int_60_141 bl_int_59_141 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c142
+ bl_int_60_142 bl_int_59_142 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c143
+ bl_int_60_143 bl_int_59_143 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c144
+ bl_int_60_144 bl_int_59_144 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c145
+ bl_int_60_145 bl_int_59_145 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c146
+ bl_int_60_146 bl_int_59_146 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c147
+ bl_int_60_147 bl_int_59_147 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c148
+ bl_int_60_148 bl_int_59_148 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c149
+ bl_int_60_149 bl_int_59_149 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c150
+ bl_int_60_150 bl_int_59_150 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c151
+ bl_int_60_151 bl_int_59_151 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c152
+ bl_int_60_152 bl_int_59_152 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c153
+ bl_int_60_153 bl_int_59_153 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c154
+ bl_int_60_154 bl_int_59_154 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c155
+ bl_int_60_155 bl_int_59_155 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c156
+ bl_int_60_156 bl_int_59_156 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c157
+ bl_int_60_157 bl_int_59_157 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c158
+ bl_int_60_158 bl_int_59_158 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c159
+ bl_int_60_159 bl_int_59_159 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c160
+ bl_int_60_160 bl_int_59_160 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c161
+ bl_int_60_161 bl_int_59_161 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c162
+ bl_int_60_162 bl_int_59_162 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c163
+ bl_int_60_163 bl_int_59_163 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c164
+ bl_int_60_164 bl_int_59_164 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c165
+ bl_int_60_165 bl_int_59_165 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c166
+ bl_int_60_166 bl_int_59_166 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c167
+ bl_int_60_167 bl_int_59_167 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c168
+ bl_int_60_168 bl_int_59_168 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c169
+ bl_int_60_169 bl_int_59_169 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c170
+ bl_int_60_170 bl_int_59_170 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c171
+ bl_int_60_171 bl_int_59_171 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c172
+ bl_int_60_172 bl_int_59_172 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c173
+ bl_int_60_173 bl_int_59_173 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c174
+ bl_int_60_174 bl_int_59_174 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c175
+ bl_int_60_175 bl_int_59_175 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c176
+ bl_int_60_176 bl_int_59_176 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c177
+ bl_int_60_177 bl_int_59_177 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c178
+ bl_int_60_178 bl_int_59_178 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c179
+ bl_int_60_179 bl_int_59_179 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c180
+ bl_int_60_180 bl_int_59_180 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c181
+ bl_int_60_181 bl_int_59_181 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c182
+ bl_int_60_182 bl_int_59_182 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r60_c183
+ bl_int_60_183 bl_int_59_183 wl_0_60 gnd
+ sram_rom_base_one_cell
Xbit_r61_c0
+ bl_int_61_0 bl_int_60_0 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c1
+ bl_int_61_1 bl_int_60_1 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c2
+ bl_int_61_2 bl_int_60_2 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c3
+ bl_int_61_3 bl_int_60_3 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c4
+ bl_int_61_4 bl_int_60_4 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c5
+ bl_int_61_5 bl_int_60_5 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c6
+ bl_int_61_6 bl_int_60_6 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c7
+ bl_int_61_7 bl_int_60_7 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c8
+ bl_int_61_8 bl_int_60_8 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c9
+ bl_int_61_9 bl_int_60_9 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c10
+ bl_int_61_10 bl_int_60_10 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c11
+ bl_int_61_11 bl_int_60_11 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c12
+ bl_int_61_12 bl_int_60_12 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c13
+ bl_int_61_13 bl_int_60_13 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c14
+ bl_int_61_14 bl_int_60_14 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c15
+ bl_int_61_15 bl_int_60_15 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c16
+ bl_int_61_16 bl_int_60_16 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c17
+ bl_int_61_17 bl_int_60_17 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c18
+ bl_int_61_18 bl_int_60_18 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c19
+ bl_int_61_19 bl_int_60_19 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c20
+ bl_int_61_20 bl_int_60_20 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c21
+ bl_int_61_21 bl_int_60_21 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c22
+ bl_int_61_22 bl_int_60_22 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c23
+ bl_int_61_23 bl_int_60_23 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c24
+ bl_int_61_24 bl_int_60_24 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c25
+ bl_int_61_25 bl_int_60_25 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c26
+ bl_int_61_26 bl_int_60_26 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c27
+ bl_int_61_27 bl_int_60_27 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c28
+ bl_int_61_28 bl_int_60_28 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c29
+ bl_int_61_29 bl_int_60_29 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c30
+ bl_int_61_30 bl_int_60_30 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c31
+ bl_int_61_31 bl_int_60_31 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c32
+ bl_int_61_32 bl_int_60_32 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c33
+ bl_int_61_33 bl_int_60_33 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c34
+ bl_int_61_34 bl_int_60_34 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c35
+ bl_int_61_35 bl_int_60_35 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c36
+ bl_int_61_36 bl_int_60_36 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c37
+ bl_int_61_37 bl_int_60_37 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c38
+ bl_int_61_38 bl_int_60_38 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c39
+ bl_int_61_39 bl_int_60_39 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c40
+ bl_int_61_40 bl_int_60_40 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c41
+ bl_int_61_41 bl_int_60_41 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c42
+ bl_int_61_42 bl_int_60_42 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c43
+ bl_int_61_43 bl_int_60_43 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c44
+ bl_int_61_44 bl_int_60_44 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c45
+ bl_int_61_45 bl_int_60_45 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c46
+ bl_int_61_46 bl_int_60_46 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c47
+ bl_int_61_47 bl_int_60_47 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c48
+ bl_int_61_48 bl_int_60_48 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c49
+ bl_int_61_49 bl_int_60_49 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c50
+ bl_int_61_50 bl_int_60_50 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c51
+ bl_int_61_51 bl_int_60_51 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c52
+ bl_int_61_52 bl_int_60_52 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c53
+ bl_int_61_53 bl_int_60_53 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c54
+ bl_int_61_54 bl_int_60_54 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c55
+ bl_int_61_55 bl_int_60_55 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c56
+ bl_int_61_56 bl_int_60_56 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c57
+ bl_int_61_57 bl_int_60_57 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c58
+ bl_int_61_58 bl_int_60_58 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c59
+ bl_int_61_59 bl_int_60_59 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c60
+ bl_int_61_60 bl_int_60_60 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c61
+ bl_int_61_61 bl_int_60_61 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c62
+ bl_int_61_62 bl_int_60_62 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c63
+ bl_int_61_63 bl_int_60_63 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c64
+ bl_int_61_64 bl_int_60_64 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c65
+ bl_int_61_65 bl_int_60_65 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c66
+ bl_int_61_66 bl_int_60_66 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c67
+ bl_int_61_67 bl_int_60_67 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c68
+ bl_int_61_68 bl_int_60_68 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c69
+ bl_int_61_69 bl_int_60_69 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c70
+ bl_int_61_70 bl_int_60_70 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c71
+ bl_int_61_71 bl_int_60_71 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c72
+ bl_int_61_72 bl_int_60_72 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c73
+ bl_int_61_73 bl_int_60_73 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c74
+ bl_int_61_74 bl_int_60_74 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c75
+ bl_int_61_75 bl_int_60_75 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c76
+ bl_int_61_76 bl_int_60_76 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c77
+ bl_int_61_77 bl_int_60_77 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c78
+ bl_int_61_78 bl_int_60_78 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c79
+ bl_int_61_79 bl_int_60_79 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c80
+ bl_int_61_80 bl_int_60_80 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c81
+ bl_int_61_81 bl_int_60_81 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c82
+ bl_int_61_82 bl_int_60_82 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c83
+ bl_int_61_83 bl_int_60_83 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c84
+ bl_int_61_84 bl_int_60_84 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c85
+ bl_int_61_85 bl_int_60_85 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c86
+ bl_int_61_86 bl_int_60_86 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c87
+ bl_int_61_87 bl_int_60_87 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c88
+ bl_int_61_88 bl_int_60_88 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c89
+ bl_int_61_89 bl_int_60_89 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c90
+ bl_int_61_90 bl_int_60_90 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c91
+ bl_int_61_91 bl_int_60_91 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c92
+ bl_int_61_92 bl_int_60_92 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c93
+ bl_int_61_93 bl_int_60_93 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c94
+ bl_int_61_94 bl_int_60_94 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c95
+ bl_int_61_95 bl_int_60_95 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c96
+ bl_int_61_96 bl_int_60_96 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c97
+ bl_int_61_97 bl_int_60_97 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c98
+ bl_int_61_98 bl_int_60_98 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c99
+ bl_int_61_99 bl_int_60_99 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c100
+ bl_int_61_100 bl_int_60_100 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c101
+ bl_int_61_101 bl_int_60_101 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c102
+ bl_int_61_102 bl_int_60_102 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c103
+ bl_int_61_103 bl_int_60_103 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c104
+ bl_int_61_104 bl_int_60_104 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c105
+ bl_int_61_105 bl_int_60_105 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c106
+ bl_int_61_106 bl_int_60_106 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c107
+ bl_int_61_107 bl_int_60_107 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c108
+ bl_int_61_108 bl_int_60_108 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c109
+ bl_int_61_109 bl_int_60_109 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c110
+ bl_int_61_110 bl_int_60_110 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c111
+ bl_int_61_111 bl_int_60_111 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c112
+ bl_int_61_112 bl_int_60_112 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c113
+ bl_int_61_113 bl_int_60_113 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c114
+ bl_int_61_114 bl_int_60_114 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c115
+ bl_int_61_115 bl_int_60_115 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c116
+ bl_int_61_116 bl_int_60_116 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c117
+ bl_int_61_117 bl_int_60_117 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c118
+ bl_int_61_118 bl_int_60_118 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c119
+ bl_int_61_119 bl_int_60_119 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c120
+ bl_int_61_120 bl_int_60_120 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c121
+ bl_int_61_121 bl_int_60_121 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c122
+ bl_int_61_122 bl_int_60_122 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c123
+ bl_int_61_123 bl_int_60_123 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c124
+ bl_int_61_124 bl_int_60_124 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c125
+ bl_int_61_125 bl_int_60_125 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c126
+ bl_int_61_126 bl_int_60_126 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c127
+ bl_int_61_127 bl_int_60_127 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c128
+ bl_int_61_128 bl_int_60_128 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c129
+ bl_int_61_129 bl_int_60_129 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c130
+ bl_int_61_130 bl_int_60_130 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c131
+ bl_int_61_131 bl_int_60_131 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c132
+ bl_int_61_132 bl_int_60_132 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c133
+ bl_int_61_133 bl_int_60_133 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c134
+ bl_int_61_134 bl_int_60_134 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c135
+ bl_int_61_135 bl_int_60_135 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c136
+ bl_int_61_136 bl_int_60_136 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c137
+ bl_int_61_137 bl_int_60_137 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c138
+ bl_int_61_138 bl_int_60_138 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c139
+ bl_int_61_139 bl_int_60_139 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c140
+ bl_int_61_140 bl_int_60_140 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c141
+ bl_int_61_141 bl_int_60_141 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c142
+ bl_int_61_142 bl_int_60_142 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c143
+ bl_int_61_143 bl_int_60_143 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c144
+ bl_int_61_144 bl_int_60_144 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c145
+ bl_int_61_145 bl_int_60_145 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c146
+ bl_int_61_146 bl_int_60_146 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c147
+ bl_int_61_147 bl_int_60_147 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c148
+ bl_int_61_148 bl_int_60_148 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c149
+ bl_int_61_149 bl_int_60_149 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c150
+ bl_int_61_150 bl_int_60_150 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c151
+ bl_int_61_151 bl_int_60_151 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c152
+ bl_int_61_152 bl_int_60_152 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c153
+ bl_int_61_153 bl_int_60_153 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c154
+ bl_int_61_154 bl_int_60_154 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c155
+ bl_int_61_155 bl_int_60_155 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c156
+ bl_int_61_156 bl_int_60_156 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c157
+ bl_int_61_157 bl_int_60_157 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c158
+ bl_int_61_158 bl_int_60_158 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c159
+ bl_int_61_159 bl_int_60_159 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c160
+ bl_int_61_160 bl_int_60_160 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c161
+ bl_int_61_161 bl_int_60_161 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c162
+ bl_int_61_162 bl_int_60_162 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c163
+ bl_int_61_163 bl_int_60_163 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c164
+ bl_int_61_164 bl_int_60_164 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c165
+ bl_int_61_165 bl_int_60_165 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c166
+ bl_int_61_166 bl_int_60_166 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c167
+ bl_int_61_167 bl_int_60_167 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c168
+ bl_int_61_168 bl_int_60_168 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c169
+ bl_int_61_169 bl_int_60_169 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c170
+ bl_int_61_170 bl_int_60_170 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c171
+ bl_int_61_171 bl_int_60_171 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c172
+ bl_int_61_172 bl_int_60_172 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c173
+ bl_int_61_173 bl_int_60_173 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c174
+ bl_int_61_174 bl_int_60_174 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c175
+ bl_int_61_175 bl_int_60_175 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c176
+ bl_int_61_176 bl_int_60_176 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c177
+ bl_int_61_177 bl_int_60_177 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c178
+ bl_int_61_178 bl_int_60_178 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c179
+ bl_int_61_179 bl_int_60_179 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c180
+ bl_int_61_180 bl_int_60_180 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c181
+ bl_int_61_181 bl_int_60_181 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c182
+ bl_int_61_182 bl_int_60_182 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r61_c183
+ bl_int_61_183 bl_int_60_183 wl_0_61 gnd
+ sram_rom_base_one_cell
Xbit_r62_c0
+ bl_int_62_0 bl_int_61_0 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c1
+ bl_int_62_1 bl_int_61_1 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c2
+ bl_int_62_2 bl_int_61_2 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c3
+ bl_int_62_3 bl_int_61_3 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c4
+ bl_int_62_4 bl_int_61_4 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c5
+ bl_int_62_5 bl_int_61_5 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c6
+ bl_int_62_6 bl_int_61_6 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c7
+ bl_int_62_7 bl_int_61_7 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c8
+ bl_int_62_8 bl_int_61_8 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c9
+ bl_int_62_9 bl_int_61_9 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c10
+ bl_int_62_10 bl_int_61_10 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c11
+ bl_int_62_11 bl_int_61_11 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c12
+ bl_int_62_12 bl_int_61_12 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c13
+ bl_int_62_13 bl_int_61_13 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c14
+ bl_int_62_14 bl_int_61_14 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c15
+ bl_int_62_15 bl_int_61_15 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c16
+ bl_int_62_16 bl_int_61_16 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c17
+ bl_int_62_17 bl_int_61_17 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c18
+ bl_int_62_18 bl_int_61_18 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c19
+ bl_int_62_19 bl_int_61_19 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c20
+ bl_int_62_20 bl_int_61_20 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c21
+ bl_int_62_21 bl_int_61_21 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c22
+ bl_int_62_22 bl_int_61_22 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c23
+ bl_int_62_23 bl_int_61_23 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c24
+ bl_int_62_24 bl_int_61_24 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c25
+ bl_int_62_25 bl_int_61_25 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c26
+ bl_int_62_26 bl_int_61_26 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c27
+ bl_int_62_27 bl_int_61_27 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c28
+ bl_int_62_28 bl_int_61_28 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c29
+ bl_int_62_29 bl_int_61_29 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c30
+ bl_int_62_30 bl_int_61_30 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c31
+ bl_int_62_31 bl_int_61_31 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c32
+ bl_int_62_32 bl_int_61_32 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c33
+ bl_int_62_33 bl_int_61_33 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c34
+ bl_int_62_34 bl_int_61_34 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c35
+ bl_int_62_35 bl_int_61_35 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c36
+ bl_int_62_36 bl_int_61_36 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c37
+ bl_int_62_37 bl_int_61_37 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c38
+ bl_int_62_38 bl_int_61_38 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c39
+ bl_int_62_39 bl_int_61_39 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c40
+ bl_int_62_40 bl_int_61_40 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c41
+ bl_int_62_41 bl_int_61_41 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c42
+ bl_int_62_42 bl_int_61_42 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c43
+ bl_int_62_43 bl_int_61_43 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c44
+ bl_int_62_44 bl_int_61_44 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c45
+ bl_int_62_45 bl_int_61_45 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c46
+ bl_int_62_46 bl_int_61_46 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c47
+ bl_int_62_47 bl_int_61_47 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c48
+ bl_int_62_48 bl_int_61_48 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c49
+ bl_int_62_49 bl_int_61_49 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c50
+ bl_int_62_50 bl_int_61_50 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c51
+ bl_int_62_51 bl_int_61_51 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c52
+ bl_int_62_52 bl_int_61_52 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c53
+ bl_int_62_53 bl_int_61_53 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c54
+ bl_int_62_54 bl_int_61_54 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c55
+ bl_int_62_55 bl_int_61_55 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c56
+ bl_int_62_56 bl_int_61_56 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c57
+ bl_int_62_57 bl_int_61_57 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c58
+ bl_int_62_58 bl_int_61_58 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c59
+ bl_int_62_59 bl_int_61_59 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c60
+ bl_int_62_60 bl_int_61_60 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c61
+ bl_int_62_61 bl_int_61_61 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c62
+ bl_int_62_62 bl_int_61_62 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c63
+ bl_int_62_63 bl_int_61_63 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c64
+ bl_int_62_64 bl_int_61_64 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c65
+ bl_int_62_65 bl_int_61_65 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c66
+ bl_int_62_66 bl_int_61_66 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c67
+ bl_int_62_67 bl_int_61_67 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c68
+ bl_int_62_68 bl_int_61_68 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c69
+ bl_int_62_69 bl_int_61_69 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c70
+ bl_int_62_70 bl_int_61_70 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c71
+ bl_int_62_71 bl_int_61_71 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c72
+ bl_int_62_72 bl_int_61_72 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c73
+ bl_int_62_73 bl_int_61_73 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c74
+ bl_int_62_74 bl_int_61_74 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c75
+ bl_int_62_75 bl_int_61_75 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c76
+ bl_int_62_76 bl_int_61_76 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c77
+ bl_int_62_77 bl_int_61_77 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c78
+ bl_int_62_78 bl_int_61_78 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c79
+ bl_int_62_79 bl_int_61_79 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c80
+ bl_int_62_80 bl_int_61_80 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c81
+ bl_int_62_81 bl_int_61_81 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c82
+ bl_int_62_82 bl_int_61_82 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c83
+ bl_int_62_83 bl_int_61_83 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c84
+ bl_int_62_84 bl_int_61_84 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c85
+ bl_int_62_85 bl_int_61_85 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c86
+ bl_int_62_86 bl_int_61_86 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c87
+ bl_int_62_87 bl_int_61_87 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c88
+ bl_int_62_88 bl_int_61_88 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c89
+ bl_int_62_89 bl_int_61_89 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c90
+ bl_int_62_90 bl_int_61_90 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c91
+ bl_int_62_91 bl_int_61_91 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c92
+ bl_int_62_92 bl_int_61_92 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c93
+ bl_int_62_93 bl_int_61_93 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c94
+ bl_int_62_94 bl_int_61_94 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c95
+ bl_int_62_95 bl_int_61_95 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c96
+ bl_int_62_96 bl_int_61_96 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c97
+ bl_int_62_97 bl_int_61_97 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c98
+ bl_int_62_98 bl_int_61_98 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c99
+ bl_int_62_99 bl_int_61_99 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c100
+ bl_int_62_100 bl_int_61_100 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c101
+ bl_int_62_101 bl_int_61_101 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c102
+ bl_int_62_102 bl_int_61_102 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c103
+ bl_int_62_103 bl_int_61_103 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c104
+ bl_int_62_104 bl_int_61_104 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c105
+ bl_int_62_105 bl_int_61_105 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c106
+ bl_int_62_106 bl_int_61_106 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c107
+ bl_int_62_107 bl_int_61_107 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c108
+ bl_int_62_108 bl_int_61_108 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c109
+ bl_int_62_109 bl_int_61_109 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c110
+ bl_int_62_110 bl_int_61_110 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c111
+ bl_int_62_111 bl_int_61_111 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c112
+ bl_int_62_112 bl_int_61_112 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c113
+ bl_int_62_113 bl_int_61_113 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c114
+ bl_int_62_114 bl_int_61_114 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c115
+ bl_int_62_115 bl_int_61_115 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c116
+ bl_int_62_116 bl_int_61_116 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c117
+ bl_int_62_117 bl_int_61_117 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c118
+ bl_int_62_118 bl_int_61_118 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c119
+ bl_int_62_119 bl_int_61_119 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c120
+ bl_int_62_120 bl_int_61_120 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c121
+ bl_int_62_121 bl_int_61_121 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c122
+ bl_int_62_122 bl_int_61_122 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c123
+ bl_int_62_123 bl_int_61_123 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c124
+ bl_int_62_124 bl_int_61_124 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c125
+ bl_int_62_125 bl_int_61_125 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c126
+ bl_int_62_126 bl_int_61_126 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c127
+ bl_int_62_127 bl_int_61_127 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c128
+ bl_int_62_128 bl_int_61_128 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c129
+ bl_int_62_129 bl_int_61_129 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c130
+ bl_int_62_130 bl_int_61_130 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c131
+ bl_int_62_131 bl_int_61_131 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c132
+ bl_int_62_132 bl_int_61_132 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c133
+ bl_int_62_133 bl_int_61_133 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c134
+ bl_int_62_134 bl_int_61_134 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c135
+ bl_int_62_135 bl_int_61_135 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c136
+ bl_int_62_136 bl_int_61_136 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c137
+ bl_int_62_137 bl_int_61_137 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c138
+ bl_int_62_138 bl_int_61_138 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c139
+ bl_int_62_139 bl_int_61_139 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c140
+ bl_int_62_140 bl_int_61_140 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c141
+ bl_int_62_141 bl_int_61_141 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c142
+ bl_int_62_142 bl_int_61_142 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c143
+ bl_int_62_143 bl_int_61_143 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c144
+ bl_int_62_144 bl_int_61_144 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c145
+ bl_int_62_145 bl_int_61_145 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c146
+ bl_int_62_146 bl_int_61_146 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c147
+ bl_int_62_147 bl_int_61_147 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c148
+ bl_int_62_148 bl_int_61_148 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c149
+ bl_int_62_149 bl_int_61_149 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c150
+ bl_int_62_150 bl_int_61_150 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c151
+ bl_int_62_151 bl_int_61_151 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c152
+ bl_int_62_152 bl_int_61_152 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c153
+ bl_int_62_153 bl_int_61_153 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c154
+ bl_int_62_154 bl_int_61_154 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c155
+ bl_int_62_155 bl_int_61_155 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c156
+ bl_int_62_156 bl_int_61_156 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c157
+ bl_int_62_157 bl_int_61_157 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c158
+ bl_int_62_158 bl_int_61_158 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c159
+ bl_int_62_159 bl_int_61_159 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c160
+ bl_int_62_160 bl_int_61_160 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c161
+ bl_int_62_161 bl_int_61_161 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c162
+ bl_int_62_162 bl_int_61_162 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c163
+ bl_int_62_163 bl_int_61_163 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c164
+ bl_int_62_164 bl_int_61_164 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c165
+ bl_int_62_165 bl_int_61_165 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c166
+ bl_int_62_166 bl_int_61_166 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c167
+ bl_int_62_167 bl_int_61_167 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c168
+ bl_int_62_168 bl_int_61_168 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c169
+ bl_int_62_169 bl_int_61_169 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c170
+ bl_int_62_170 bl_int_61_170 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c171
+ bl_int_62_171 bl_int_61_171 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c172
+ bl_int_62_172 bl_int_61_172 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c173
+ bl_int_62_173 bl_int_61_173 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c174
+ bl_int_62_174 bl_int_61_174 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c175
+ bl_int_62_175 bl_int_61_175 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c176
+ bl_int_62_176 bl_int_61_176 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c177
+ bl_int_62_177 bl_int_61_177 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c178
+ bl_int_62_178 bl_int_61_178 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c179
+ bl_int_62_179 bl_int_61_179 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c180
+ bl_int_62_180 bl_int_61_180 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c181
+ bl_int_62_181 bl_int_61_181 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c182
+ bl_int_62_182 bl_int_61_182 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r62_c183
+ bl_int_62_183 bl_int_61_183 wl_0_62 gnd
+ sram_rom_base_one_cell
Xbit_r63_c0
+ bl_int_63_0 bl_int_62_0 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c1
+ bl_int_63_1 bl_int_62_1 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c2
+ bl_int_63_2 bl_int_62_2 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c3
+ bl_int_63_3 bl_int_62_3 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c4
+ bl_int_63_4 bl_int_62_4 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c5
+ bl_int_63_5 bl_int_62_5 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c6
+ bl_int_63_6 bl_int_62_6 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c7
+ bl_int_63_7 bl_int_62_7 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c8
+ bl_int_63_8 bl_int_62_8 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c9
+ bl_int_63_9 bl_int_62_9 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c10
+ bl_int_63_10 bl_int_62_10 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c11
+ bl_int_63_11 bl_int_62_11 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c12
+ bl_int_63_12 bl_int_62_12 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c13
+ bl_int_63_13 bl_int_62_13 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c14
+ bl_int_63_14 bl_int_62_14 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c15
+ bl_int_63_15 bl_int_62_15 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c16
+ bl_int_63_16 bl_int_62_16 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c17
+ bl_int_63_17 bl_int_62_17 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c18
+ bl_int_63_18 bl_int_62_18 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c19
+ bl_int_63_19 bl_int_62_19 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c20
+ bl_int_63_20 bl_int_62_20 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c21
+ bl_int_63_21 bl_int_62_21 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c22
+ bl_int_63_22 bl_int_62_22 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c23
+ bl_int_63_23 bl_int_62_23 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c24
+ bl_int_63_24 bl_int_62_24 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c25
+ bl_int_63_25 bl_int_62_25 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c26
+ bl_int_63_26 bl_int_62_26 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c27
+ bl_int_63_27 bl_int_62_27 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c28
+ bl_int_63_28 bl_int_62_28 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c29
+ bl_int_63_29 bl_int_62_29 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c30
+ bl_int_63_30 bl_int_62_30 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c31
+ bl_int_63_31 bl_int_62_31 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c32
+ bl_int_63_32 bl_int_62_32 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c33
+ bl_int_63_33 bl_int_62_33 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c34
+ bl_int_63_34 bl_int_62_34 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c35
+ bl_int_63_35 bl_int_62_35 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c36
+ bl_int_63_36 bl_int_62_36 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c37
+ bl_int_63_37 bl_int_62_37 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c38
+ bl_int_63_38 bl_int_62_38 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c39
+ bl_int_63_39 bl_int_62_39 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c40
+ bl_int_63_40 bl_int_62_40 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c41
+ bl_int_63_41 bl_int_62_41 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c42
+ bl_int_63_42 bl_int_62_42 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c43
+ bl_int_63_43 bl_int_62_43 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c44
+ bl_int_63_44 bl_int_62_44 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c45
+ bl_int_63_45 bl_int_62_45 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c46
+ bl_int_63_46 bl_int_62_46 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c47
+ bl_int_63_47 bl_int_62_47 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c48
+ bl_int_63_48 bl_int_62_48 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c49
+ bl_int_63_49 bl_int_62_49 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c50
+ bl_int_63_50 bl_int_62_50 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c51
+ bl_int_63_51 bl_int_62_51 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c52
+ bl_int_63_52 bl_int_62_52 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c53
+ bl_int_63_53 bl_int_62_53 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c54
+ bl_int_63_54 bl_int_62_54 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c55
+ bl_int_63_55 bl_int_62_55 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c56
+ bl_int_63_56 bl_int_62_56 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c57
+ bl_int_63_57 bl_int_62_57 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c58
+ bl_int_63_58 bl_int_62_58 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c59
+ bl_int_63_59 bl_int_62_59 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c60
+ bl_int_63_60 bl_int_62_60 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c61
+ bl_int_63_61 bl_int_62_61 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c62
+ bl_int_63_62 bl_int_62_62 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c63
+ bl_int_63_63 bl_int_62_63 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c64
+ bl_int_63_64 bl_int_62_64 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c65
+ bl_int_63_65 bl_int_62_65 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c66
+ bl_int_63_66 bl_int_62_66 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c67
+ bl_int_63_67 bl_int_62_67 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c68
+ bl_int_63_68 bl_int_62_68 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c69
+ bl_int_63_69 bl_int_62_69 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c70
+ bl_int_63_70 bl_int_62_70 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c71
+ bl_int_63_71 bl_int_62_71 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c72
+ bl_int_63_72 bl_int_62_72 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c73
+ bl_int_63_73 bl_int_62_73 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c74
+ bl_int_63_74 bl_int_62_74 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c75
+ bl_int_63_75 bl_int_62_75 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c76
+ bl_int_63_76 bl_int_62_76 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c77
+ bl_int_63_77 bl_int_62_77 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c78
+ bl_int_63_78 bl_int_62_78 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c79
+ bl_int_63_79 bl_int_62_79 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c80
+ bl_int_63_80 bl_int_62_80 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c81
+ bl_int_63_81 bl_int_62_81 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c82
+ bl_int_63_82 bl_int_62_82 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c83
+ bl_int_63_83 bl_int_62_83 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c84
+ bl_int_63_84 bl_int_62_84 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c85
+ bl_int_63_85 bl_int_62_85 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c86
+ bl_int_63_86 bl_int_62_86 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c87
+ bl_int_63_87 bl_int_62_87 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c88
+ bl_int_63_88 bl_int_62_88 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c89
+ bl_int_63_89 bl_int_62_89 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c90
+ bl_int_63_90 bl_int_62_90 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c91
+ bl_int_63_91 bl_int_62_91 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c92
+ bl_int_63_92 bl_int_62_92 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c93
+ bl_int_63_93 bl_int_62_93 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c94
+ bl_int_63_94 bl_int_62_94 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c95
+ bl_int_63_95 bl_int_62_95 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c96
+ bl_int_63_96 bl_int_62_96 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c97
+ bl_int_63_97 bl_int_62_97 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c98
+ bl_int_63_98 bl_int_62_98 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c99
+ bl_int_63_99 bl_int_62_99 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c100
+ bl_int_63_100 bl_int_62_100 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c101
+ bl_int_63_101 bl_int_62_101 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c102
+ bl_int_63_102 bl_int_62_102 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c103
+ bl_int_63_103 bl_int_62_103 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c104
+ bl_int_63_104 bl_int_62_104 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c105
+ bl_int_63_105 bl_int_62_105 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c106
+ bl_int_63_106 bl_int_62_106 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c107
+ bl_int_63_107 bl_int_62_107 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c108
+ bl_int_63_108 bl_int_62_108 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c109
+ bl_int_63_109 bl_int_62_109 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c110
+ bl_int_63_110 bl_int_62_110 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c111
+ bl_int_63_111 bl_int_62_111 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c112
+ bl_int_63_112 bl_int_62_112 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c113
+ bl_int_63_113 bl_int_62_113 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c114
+ bl_int_63_114 bl_int_62_114 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c115
+ bl_int_63_115 bl_int_62_115 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c116
+ bl_int_63_116 bl_int_62_116 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c117
+ bl_int_63_117 bl_int_62_117 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c118
+ bl_int_63_118 bl_int_62_118 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c119
+ bl_int_63_119 bl_int_62_119 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c120
+ bl_int_63_120 bl_int_62_120 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c121
+ bl_int_63_121 bl_int_62_121 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c122
+ bl_int_63_122 bl_int_62_122 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c123
+ bl_int_63_123 bl_int_62_123 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c124
+ bl_int_63_124 bl_int_62_124 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c125
+ bl_int_63_125 bl_int_62_125 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c126
+ bl_int_63_126 bl_int_62_126 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c127
+ bl_int_63_127 bl_int_62_127 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c128
+ bl_int_63_128 bl_int_62_128 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c129
+ bl_int_63_129 bl_int_62_129 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c130
+ bl_int_63_130 bl_int_62_130 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c131
+ bl_int_63_131 bl_int_62_131 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c132
+ bl_int_63_132 bl_int_62_132 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c133
+ bl_int_63_133 bl_int_62_133 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c134
+ bl_int_63_134 bl_int_62_134 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c135
+ bl_int_63_135 bl_int_62_135 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c136
+ bl_int_63_136 bl_int_62_136 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c137
+ bl_int_63_137 bl_int_62_137 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c138
+ bl_int_63_138 bl_int_62_138 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c139
+ bl_int_63_139 bl_int_62_139 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c140
+ bl_int_63_140 bl_int_62_140 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c141
+ bl_int_63_141 bl_int_62_141 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c142
+ bl_int_63_142 bl_int_62_142 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c143
+ bl_int_63_143 bl_int_62_143 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c144
+ bl_int_63_144 bl_int_62_144 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c145
+ bl_int_63_145 bl_int_62_145 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c146
+ bl_int_63_146 bl_int_62_146 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c147
+ bl_int_63_147 bl_int_62_147 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c148
+ bl_int_63_148 bl_int_62_148 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c149
+ bl_int_63_149 bl_int_62_149 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c150
+ bl_int_63_150 bl_int_62_150 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c151
+ bl_int_63_151 bl_int_62_151 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c152
+ bl_int_63_152 bl_int_62_152 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c153
+ bl_int_63_153 bl_int_62_153 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c154
+ bl_int_63_154 bl_int_62_154 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c155
+ bl_int_63_155 bl_int_62_155 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c156
+ bl_int_63_156 bl_int_62_156 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c157
+ bl_int_63_157 bl_int_62_157 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c158
+ bl_int_63_158 bl_int_62_158 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c159
+ bl_int_63_159 bl_int_62_159 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c160
+ bl_int_63_160 bl_int_62_160 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c161
+ bl_int_63_161 bl_int_62_161 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c162
+ bl_int_63_162 bl_int_62_162 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c163
+ bl_int_63_163 bl_int_62_163 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c164
+ bl_int_63_164 bl_int_62_164 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c165
+ bl_int_63_165 bl_int_62_165 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c166
+ bl_int_63_166 bl_int_62_166 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c167
+ bl_int_63_167 bl_int_62_167 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c168
+ bl_int_63_168 bl_int_62_168 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c169
+ bl_int_63_169 bl_int_62_169 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c170
+ bl_int_63_170 bl_int_62_170 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c171
+ bl_int_63_171 bl_int_62_171 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c172
+ bl_int_63_172 bl_int_62_172 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c173
+ bl_int_63_173 bl_int_62_173 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c174
+ bl_int_63_174 bl_int_62_174 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c175
+ bl_int_63_175 bl_int_62_175 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c176
+ bl_int_63_176 bl_int_62_176 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c177
+ bl_int_63_177 bl_int_62_177 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c178
+ bl_int_63_178 bl_int_62_178 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c179
+ bl_int_63_179 bl_int_62_179 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c180
+ bl_int_63_180 bl_int_62_180 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c181
+ bl_int_63_181 bl_int_62_181 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c182
+ bl_int_63_182 bl_int_62_182 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r63_c183
+ bl_int_63_183 bl_int_62_183 wl_0_63 gnd
+ sram_rom_base_one_cell
Xbit_r64_c0
+ bl_int_64_0 bl_int_63_0 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c1
+ bl_int_64_1 bl_int_63_1 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c2
+ bl_int_64_2 bl_int_63_2 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c3
+ bl_int_64_3 bl_int_63_3 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c4
+ bl_int_64_4 bl_int_63_4 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c5
+ bl_int_64_5 bl_int_63_5 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c6
+ bl_int_64_6 bl_int_63_6 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c7
+ bl_int_64_7 bl_int_63_7 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c8
+ bl_int_64_8 bl_int_63_8 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c9
+ bl_int_64_9 bl_int_63_9 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c10
+ bl_int_64_10 bl_int_63_10 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c11
+ bl_int_64_11 bl_int_63_11 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c12
+ bl_int_64_12 bl_int_63_12 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c13
+ bl_int_64_13 bl_int_63_13 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c14
+ bl_int_64_14 bl_int_63_14 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c15
+ bl_int_64_15 bl_int_63_15 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c16
+ bl_int_64_16 bl_int_63_16 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c17
+ bl_int_64_17 bl_int_63_17 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c18
+ bl_int_64_18 bl_int_63_18 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c19
+ bl_int_64_19 bl_int_63_19 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c20
+ bl_int_64_20 bl_int_63_20 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c21
+ bl_int_64_21 bl_int_63_21 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c22
+ bl_int_64_22 bl_int_63_22 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c23
+ bl_int_64_23 bl_int_63_23 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c24
+ bl_int_64_24 bl_int_63_24 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c25
+ bl_int_64_25 bl_int_63_25 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c26
+ bl_int_64_26 bl_int_63_26 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c27
+ bl_int_64_27 bl_int_63_27 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c28
+ bl_int_64_28 bl_int_63_28 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c29
+ bl_int_64_29 bl_int_63_29 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c30
+ bl_int_64_30 bl_int_63_30 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c31
+ bl_int_64_31 bl_int_63_31 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c32
+ bl_int_64_32 bl_int_63_32 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c33
+ bl_int_64_33 bl_int_63_33 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c34
+ bl_int_64_34 bl_int_63_34 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c35
+ bl_int_64_35 bl_int_63_35 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c36
+ bl_int_64_36 bl_int_63_36 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c37
+ bl_int_64_37 bl_int_63_37 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c38
+ bl_int_64_38 bl_int_63_38 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c39
+ bl_int_64_39 bl_int_63_39 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c40
+ bl_int_64_40 bl_int_63_40 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c41
+ bl_int_64_41 bl_int_63_41 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c42
+ bl_int_64_42 bl_int_63_42 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c43
+ bl_int_64_43 bl_int_63_43 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c44
+ bl_int_64_44 bl_int_63_44 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c45
+ bl_int_64_45 bl_int_63_45 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c46
+ bl_int_64_46 bl_int_63_46 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c47
+ bl_int_64_47 bl_int_63_47 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c48
+ bl_int_64_48 bl_int_63_48 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c49
+ bl_int_64_49 bl_int_63_49 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c50
+ bl_int_64_50 bl_int_63_50 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c51
+ bl_int_64_51 bl_int_63_51 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c52
+ bl_int_64_52 bl_int_63_52 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c53
+ bl_int_64_53 bl_int_63_53 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c54
+ bl_int_64_54 bl_int_63_54 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c55
+ bl_int_64_55 bl_int_63_55 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c56
+ bl_int_64_56 bl_int_63_56 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c57
+ bl_int_64_57 bl_int_63_57 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c58
+ bl_int_64_58 bl_int_63_58 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c59
+ bl_int_64_59 bl_int_63_59 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c60
+ bl_int_64_60 bl_int_63_60 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c61
+ bl_int_64_61 bl_int_63_61 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c62
+ bl_int_64_62 bl_int_63_62 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c63
+ bl_int_64_63 bl_int_63_63 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c64
+ bl_int_64_64 bl_int_63_64 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c65
+ bl_int_64_65 bl_int_63_65 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c66
+ bl_int_64_66 bl_int_63_66 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c67
+ bl_int_64_67 bl_int_63_67 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c68
+ bl_int_64_68 bl_int_63_68 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c69
+ bl_int_64_69 bl_int_63_69 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c70
+ bl_int_64_70 bl_int_63_70 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c71
+ bl_int_64_71 bl_int_63_71 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c72
+ bl_int_64_72 bl_int_63_72 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c73
+ bl_int_64_73 bl_int_63_73 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c74
+ bl_int_64_74 bl_int_63_74 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c75
+ bl_int_64_75 bl_int_63_75 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c76
+ bl_int_64_76 bl_int_63_76 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c77
+ bl_int_64_77 bl_int_63_77 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c78
+ bl_int_64_78 bl_int_63_78 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c79
+ bl_int_64_79 bl_int_63_79 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c80
+ bl_int_64_80 bl_int_63_80 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c81
+ bl_int_64_81 bl_int_63_81 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c82
+ bl_int_64_82 bl_int_63_82 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c83
+ bl_int_64_83 bl_int_63_83 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c84
+ bl_int_64_84 bl_int_63_84 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c85
+ bl_int_64_85 bl_int_63_85 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c86
+ bl_int_64_86 bl_int_63_86 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c87
+ bl_int_64_87 bl_int_63_87 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c88
+ bl_int_64_88 bl_int_63_88 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c89
+ bl_int_64_89 bl_int_63_89 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c90
+ bl_int_64_90 bl_int_63_90 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c91
+ bl_int_64_91 bl_int_63_91 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c92
+ bl_int_64_92 bl_int_63_92 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c93
+ bl_int_64_93 bl_int_63_93 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c94
+ bl_int_64_94 bl_int_63_94 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c95
+ bl_int_64_95 bl_int_63_95 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c96
+ bl_int_64_96 bl_int_63_96 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c97
+ bl_int_64_97 bl_int_63_97 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c98
+ bl_int_64_98 bl_int_63_98 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c99
+ bl_int_64_99 bl_int_63_99 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c100
+ bl_int_64_100 bl_int_63_100 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c101
+ bl_int_64_101 bl_int_63_101 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c102
+ bl_int_64_102 bl_int_63_102 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c103
+ bl_int_64_103 bl_int_63_103 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c104
+ bl_int_64_104 bl_int_63_104 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c105
+ bl_int_64_105 bl_int_63_105 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c106
+ bl_int_64_106 bl_int_63_106 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c107
+ bl_int_64_107 bl_int_63_107 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c108
+ bl_int_64_108 bl_int_63_108 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c109
+ bl_int_64_109 bl_int_63_109 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c110
+ bl_int_64_110 bl_int_63_110 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c111
+ bl_int_64_111 bl_int_63_111 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c112
+ bl_int_64_112 bl_int_63_112 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c113
+ bl_int_64_113 bl_int_63_113 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c114
+ bl_int_64_114 bl_int_63_114 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c115
+ bl_int_64_115 bl_int_63_115 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c116
+ bl_int_64_116 bl_int_63_116 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c117
+ bl_int_64_117 bl_int_63_117 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c118
+ bl_int_64_118 bl_int_63_118 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c119
+ bl_int_64_119 bl_int_63_119 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c120
+ bl_int_64_120 bl_int_63_120 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c121
+ bl_int_64_121 bl_int_63_121 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c122
+ bl_int_64_122 bl_int_63_122 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c123
+ bl_int_64_123 bl_int_63_123 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c124
+ bl_int_64_124 bl_int_63_124 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c125
+ bl_int_64_125 bl_int_63_125 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c126
+ bl_int_64_126 bl_int_63_126 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c127
+ bl_int_64_127 bl_int_63_127 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c128
+ bl_int_64_128 bl_int_63_128 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c129
+ bl_int_64_129 bl_int_63_129 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c130
+ bl_int_64_130 bl_int_63_130 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c131
+ bl_int_64_131 bl_int_63_131 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c132
+ bl_int_64_132 bl_int_63_132 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c133
+ bl_int_64_133 bl_int_63_133 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c134
+ bl_int_64_134 bl_int_63_134 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c135
+ bl_int_64_135 bl_int_63_135 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c136
+ bl_int_64_136 bl_int_63_136 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c137
+ bl_int_64_137 bl_int_63_137 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c138
+ bl_int_64_138 bl_int_63_138 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c139
+ bl_int_64_139 bl_int_63_139 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c140
+ bl_int_64_140 bl_int_63_140 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c141
+ bl_int_64_141 bl_int_63_141 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c142
+ bl_int_64_142 bl_int_63_142 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c143
+ bl_int_64_143 bl_int_63_143 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c144
+ bl_int_64_144 bl_int_63_144 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c145
+ bl_int_64_145 bl_int_63_145 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c146
+ bl_int_64_146 bl_int_63_146 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c147
+ bl_int_64_147 bl_int_63_147 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c148
+ bl_int_64_148 bl_int_63_148 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c149
+ bl_int_64_149 bl_int_63_149 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c150
+ bl_int_64_150 bl_int_63_150 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c151
+ bl_int_64_151 bl_int_63_151 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c152
+ bl_int_64_152 bl_int_63_152 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c153
+ bl_int_64_153 bl_int_63_153 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c154
+ bl_int_64_154 bl_int_63_154 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c155
+ bl_int_64_155 bl_int_63_155 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c156
+ bl_int_64_156 bl_int_63_156 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c157
+ bl_int_64_157 bl_int_63_157 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c158
+ bl_int_64_158 bl_int_63_158 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c159
+ bl_int_64_159 bl_int_63_159 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c160
+ bl_int_64_160 bl_int_63_160 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c161
+ bl_int_64_161 bl_int_63_161 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c162
+ bl_int_64_162 bl_int_63_162 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c163
+ bl_int_64_163 bl_int_63_163 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c164
+ bl_int_64_164 bl_int_63_164 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c165
+ bl_int_64_165 bl_int_63_165 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c166
+ bl_int_64_166 bl_int_63_166 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c167
+ bl_int_64_167 bl_int_63_167 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c168
+ bl_int_64_168 bl_int_63_168 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c169
+ bl_int_64_169 bl_int_63_169 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c170
+ bl_int_64_170 bl_int_63_170 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c171
+ bl_int_64_171 bl_int_63_171 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c172
+ bl_int_64_172 bl_int_63_172 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c173
+ bl_int_64_173 bl_int_63_173 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c174
+ bl_int_64_174 bl_int_63_174 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c175
+ bl_int_64_175 bl_int_63_175 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c176
+ bl_int_64_176 bl_int_63_176 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c177
+ bl_int_64_177 bl_int_63_177 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c178
+ bl_int_64_178 bl_int_63_178 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c179
+ bl_int_64_179 bl_int_63_179 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c180
+ bl_int_64_180 bl_int_63_180 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c181
+ bl_int_64_181 bl_int_63_181 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c182
+ bl_int_64_182 bl_int_63_182 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r64_c183
+ bl_int_64_183 bl_int_63_183 wl_0_64 gnd
+ sram_rom_base_one_cell
Xbit_r65_c0
+ bl_int_65_0 bl_int_64_0 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c1
+ bl_int_65_1 bl_int_64_1 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c2
+ bl_int_65_2 bl_int_64_2 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c3
+ bl_int_65_3 bl_int_64_3 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c4
+ bl_int_65_4 bl_int_64_4 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c5
+ bl_int_65_5 bl_int_64_5 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c6
+ bl_int_65_6 bl_int_64_6 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c7
+ bl_int_65_7 bl_int_64_7 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c8
+ bl_int_65_8 bl_int_64_8 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c9
+ bl_int_65_9 bl_int_64_9 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c10
+ bl_int_65_10 bl_int_64_10 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c11
+ bl_int_65_11 bl_int_64_11 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c12
+ bl_int_65_12 bl_int_64_12 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c13
+ bl_int_65_13 bl_int_64_13 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c14
+ bl_int_65_14 bl_int_64_14 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c15
+ bl_int_65_15 bl_int_64_15 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c16
+ bl_int_65_16 bl_int_64_16 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c17
+ bl_int_65_17 bl_int_64_17 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c18
+ bl_int_65_18 bl_int_64_18 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c19
+ bl_int_65_19 bl_int_64_19 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c20
+ bl_int_65_20 bl_int_64_20 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c21
+ bl_int_65_21 bl_int_64_21 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c22
+ bl_int_65_22 bl_int_64_22 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c23
+ bl_int_65_23 bl_int_64_23 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c24
+ bl_int_65_24 bl_int_64_24 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c25
+ bl_int_65_25 bl_int_64_25 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c26
+ bl_int_65_26 bl_int_64_26 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c27
+ bl_int_65_27 bl_int_64_27 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c28
+ bl_int_65_28 bl_int_64_28 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c29
+ bl_int_65_29 bl_int_64_29 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c30
+ bl_int_65_30 bl_int_64_30 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c31
+ bl_int_65_31 bl_int_64_31 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c32
+ bl_int_65_32 bl_int_64_32 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c33
+ bl_int_65_33 bl_int_64_33 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c34
+ bl_int_65_34 bl_int_64_34 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c35
+ bl_int_65_35 bl_int_64_35 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c36
+ bl_int_65_36 bl_int_64_36 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c37
+ bl_int_65_37 bl_int_64_37 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c38
+ bl_int_65_38 bl_int_64_38 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c39
+ bl_int_65_39 bl_int_64_39 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c40
+ bl_int_65_40 bl_int_64_40 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c41
+ bl_int_65_41 bl_int_64_41 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c42
+ bl_int_65_42 bl_int_64_42 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c43
+ bl_int_65_43 bl_int_64_43 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c44
+ bl_int_65_44 bl_int_64_44 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c45
+ bl_int_65_45 bl_int_64_45 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c46
+ bl_int_65_46 bl_int_64_46 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c47
+ bl_int_65_47 bl_int_64_47 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c48
+ bl_int_65_48 bl_int_64_48 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c49
+ bl_int_65_49 bl_int_64_49 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c50
+ bl_int_65_50 bl_int_64_50 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c51
+ bl_int_65_51 bl_int_64_51 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c52
+ bl_int_65_52 bl_int_64_52 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c53
+ bl_int_65_53 bl_int_64_53 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c54
+ bl_int_65_54 bl_int_64_54 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c55
+ bl_int_65_55 bl_int_64_55 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c56
+ bl_int_65_56 bl_int_64_56 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c57
+ bl_int_65_57 bl_int_64_57 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c58
+ bl_int_65_58 bl_int_64_58 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c59
+ bl_int_65_59 bl_int_64_59 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c60
+ bl_int_65_60 bl_int_64_60 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c61
+ bl_int_65_61 bl_int_64_61 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c62
+ bl_int_65_62 bl_int_64_62 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c63
+ bl_int_65_63 bl_int_64_63 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c64
+ bl_int_65_64 bl_int_64_64 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c65
+ bl_int_65_65 bl_int_64_65 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c66
+ bl_int_65_66 bl_int_64_66 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c67
+ bl_int_65_67 bl_int_64_67 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c68
+ bl_int_65_68 bl_int_64_68 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c69
+ bl_int_65_69 bl_int_64_69 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c70
+ bl_int_65_70 bl_int_64_70 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c71
+ bl_int_65_71 bl_int_64_71 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c72
+ bl_int_65_72 bl_int_64_72 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c73
+ bl_int_65_73 bl_int_64_73 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c74
+ bl_int_65_74 bl_int_64_74 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c75
+ bl_int_65_75 bl_int_64_75 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c76
+ bl_int_65_76 bl_int_64_76 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c77
+ bl_int_65_77 bl_int_64_77 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c78
+ bl_int_65_78 bl_int_64_78 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c79
+ bl_int_65_79 bl_int_64_79 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c80
+ bl_int_65_80 bl_int_64_80 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c81
+ bl_int_65_81 bl_int_64_81 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c82
+ bl_int_65_82 bl_int_64_82 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c83
+ bl_int_65_83 bl_int_64_83 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c84
+ bl_int_65_84 bl_int_64_84 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c85
+ bl_int_65_85 bl_int_64_85 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c86
+ bl_int_65_86 bl_int_64_86 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c87
+ bl_int_65_87 bl_int_64_87 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c88
+ bl_int_65_88 bl_int_64_88 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c89
+ bl_int_65_89 bl_int_64_89 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c90
+ bl_int_65_90 bl_int_64_90 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c91
+ bl_int_65_91 bl_int_64_91 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c92
+ bl_int_65_92 bl_int_64_92 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c93
+ bl_int_65_93 bl_int_64_93 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c94
+ bl_int_65_94 bl_int_64_94 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c95
+ bl_int_65_95 bl_int_64_95 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c96
+ bl_int_65_96 bl_int_64_96 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c97
+ bl_int_65_97 bl_int_64_97 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c98
+ bl_int_65_98 bl_int_64_98 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c99
+ bl_int_65_99 bl_int_64_99 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c100
+ bl_int_65_100 bl_int_64_100 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c101
+ bl_int_65_101 bl_int_64_101 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c102
+ bl_int_65_102 bl_int_64_102 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c103
+ bl_int_65_103 bl_int_64_103 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c104
+ bl_int_65_104 bl_int_64_104 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c105
+ bl_int_65_105 bl_int_64_105 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c106
+ bl_int_65_106 bl_int_64_106 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c107
+ bl_int_65_107 bl_int_64_107 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c108
+ bl_int_65_108 bl_int_64_108 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c109
+ bl_int_65_109 bl_int_64_109 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c110
+ bl_int_65_110 bl_int_64_110 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c111
+ bl_int_65_111 bl_int_64_111 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c112
+ bl_int_65_112 bl_int_64_112 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c113
+ bl_int_65_113 bl_int_64_113 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c114
+ bl_int_65_114 bl_int_64_114 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c115
+ bl_int_65_115 bl_int_64_115 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c116
+ bl_int_65_116 bl_int_64_116 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c117
+ bl_int_65_117 bl_int_64_117 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c118
+ bl_int_65_118 bl_int_64_118 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c119
+ bl_int_65_119 bl_int_64_119 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c120
+ bl_int_65_120 bl_int_64_120 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c121
+ bl_int_65_121 bl_int_64_121 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c122
+ bl_int_65_122 bl_int_64_122 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c123
+ bl_int_65_123 bl_int_64_123 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c124
+ bl_int_65_124 bl_int_64_124 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c125
+ bl_int_65_125 bl_int_64_125 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c126
+ bl_int_65_126 bl_int_64_126 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c127
+ bl_int_65_127 bl_int_64_127 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c128
+ bl_int_65_128 bl_int_64_128 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c129
+ bl_int_65_129 bl_int_64_129 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c130
+ bl_int_65_130 bl_int_64_130 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c131
+ bl_int_65_131 bl_int_64_131 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c132
+ bl_int_65_132 bl_int_64_132 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c133
+ bl_int_65_133 bl_int_64_133 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c134
+ bl_int_65_134 bl_int_64_134 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c135
+ bl_int_65_135 bl_int_64_135 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c136
+ bl_int_65_136 bl_int_64_136 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c137
+ bl_int_65_137 bl_int_64_137 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c138
+ bl_int_65_138 bl_int_64_138 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c139
+ bl_int_65_139 bl_int_64_139 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c140
+ bl_int_65_140 bl_int_64_140 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c141
+ bl_int_65_141 bl_int_64_141 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c142
+ bl_int_65_142 bl_int_64_142 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c143
+ bl_int_65_143 bl_int_64_143 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c144
+ bl_int_65_144 bl_int_64_144 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c145
+ bl_int_65_145 bl_int_64_145 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c146
+ bl_int_65_146 bl_int_64_146 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c147
+ bl_int_65_147 bl_int_64_147 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c148
+ bl_int_65_148 bl_int_64_148 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c149
+ bl_int_65_149 bl_int_64_149 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c150
+ bl_int_65_150 bl_int_64_150 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c151
+ bl_int_65_151 bl_int_64_151 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c152
+ bl_int_65_152 bl_int_64_152 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c153
+ bl_int_65_153 bl_int_64_153 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c154
+ bl_int_65_154 bl_int_64_154 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c155
+ bl_int_65_155 bl_int_64_155 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c156
+ bl_int_65_156 bl_int_64_156 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c157
+ bl_int_65_157 bl_int_64_157 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c158
+ bl_int_65_158 bl_int_64_158 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c159
+ bl_int_65_159 bl_int_64_159 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c160
+ bl_int_65_160 bl_int_64_160 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c161
+ bl_int_65_161 bl_int_64_161 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c162
+ bl_int_65_162 bl_int_64_162 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c163
+ bl_int_65_163 bl_int_64_163 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c164
+ bl_int_65_164 bl_int_64_164 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c165
+ bl_int_65_165 bl_int_64_165 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c166
+ bl_int_65_166 bl_int_64_166 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c167
+ bl_int_65_167 bl_int_64_167 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c168
+ bl_int_65_168 bl_int_64_168 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c169
+ bl_int_65_169 bl_int_64_169 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c170
+ bl_int_65_170 bl_int_64_170 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c171
+ bl_int_65_171 bl_int_64_171 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c172
+ bl_int_65_172 bl_int_64_172 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c173
+ bl_int_65_173 bl_int_64_173 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c174
+ bl_int_65_174 bl_int_64_174 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c175
+ bl_int_65_175 bl_int_64_175 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c176
+ bl_int_65_176 bl_int_64_176 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c177
+ bl_int_65_177 bl_int_64_177 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c178
+ bl_int_65_178 bl_int_64_178 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c179
+ bl_int_65_179 bl_int_64_179 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c180
+ bl_int_65_180 bl_int_64_180 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c181
+ bl_int_65_181 bl_int_64_181 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c182
+ bl_int_65_182 bl_int_64_182 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r65_c183
+ bl_int_65_183 bl_int_64_183 wl_0_65 gnd
+ sram_rom_base_one_cell
Xbit_r66_c0
+ bl_int_66_0 bl_int_65_0 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c1
+ bl_int_66_1 bl_int_65_1 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c2
+ bl_int_66_2 bl_int_65_2 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c3
+ bl_int_66_3 bl_int_65_3 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c4
+ bl_int_66_4 bl_int_65_4 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c5
+ bl_int_66_5 bl_int_65_5 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c6
+ bl_int_66_6 bl_int_65_6 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c7
+ bl_int_66_7 bl_int_65_7 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c8
+ bl_int_66_8 bl_int_65_8 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c9
+ bl_int_66_9 bl_int_65_9 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c10
+ bl_int_66_10 bl_int_65_10 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c11
+ bl_int_66_11 bl_int_65_11 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c12
+ bl_int_66_12 bl_int_65_12 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c13
+ bl_int_66_13 bl_int_65_13 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c14
+ bl_int_66_14 bl_int_65_14 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c15
+ bl_int_66_15 bl_int_65_15 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c16
+ bl_int_66_16 bl_int_65_16 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c17
+ bl_int_66_17 bl_int_65_17 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c18
+ bl_int_66_18 bl_int_65_18 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c19
+ bl_int_66_19 bl_int_65_19 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c20
+ bl_int_66_20 bl_int_65_20 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c21
+ bl_int_66_21 bl_int_65_21 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c22
+ bl_int_66_22 bl_int_65_22 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c23
+ bl_int_66_23 bl_int_65_23 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c24
+ bl_int_66_24 bl_int_65_24 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c25
+ bl_int_66_25 bl_int_65_25 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c26
+ bl_int_66_26 bl_int_65_26 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c27
+ bl_int_66_27 bl_int_65_27 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c28
+ bl_int_66_28 bl_int_65_28 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c29
+ bl_int_66_29 bl_int_65_29 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c30
+ bl_int_66_30 bl_int_65_30 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c31
+ bl_int_66_31 bl_int_65_31 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c32
+ bl_int_66_32 bl_int_65_32 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c33
+ bl_int_66_33 bl_int_65_33 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c34
+ bl_int_66_34 bl_int_65_34 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c35
+ bl_int_66_35 bl_int_65_35 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c36
+ bl_int_66_36 bl_int_65_36 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c37
+ bl_int_66_37 bl_int_65_37 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c38
+ bl_int_66_38 bl_int_65_38 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c39
+ bl_int_66_39 bl_int_65_39 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c40
+ bl_int_66_40 bl_int_65_40 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c41
+ bl_int_66_41 bl_int_65_41 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c42
+ bl_int_66_42 bl_int_65_42 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c43
+ bl_int_66_43 bl_int_65_43 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c44
+ bl_int_66_44 bl_int_65_44 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c45
+ bl_int_66_45 bl_int_65_45 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c46
+ bl_int_66_46 bl_int_65_46 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c47
+ bl_int_66_47 bl_int_65_47 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c48
+ bl_int_66_48 bl_int_65_48 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c49
+ bl_int_66_49 bl_int_65_49 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c50
+ bl_int_66_50 bl_int_65_50 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c51
+ bl_int_66_51 bl_int_65_51 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c52
+ bl_int_66_52 bl_int_65_52 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c53
+ bl_int_66_53 bl_int_65_53 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c54
+ bl_int_66_54 bl_int_65_54 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c55
+ bl_int_66_55 bl_int_65_55 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c56
+ bl_int_66_56 bl_int_65_56 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c57
+ bl_int_66_57 bl_int_65_57 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c58
+ bl_int_66_58 bl_int_65_58 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c59
+ bl_int_66_59 bl_int_65_59 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c60
+ bl_int_66_60 bl_int_65_60 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c61
+ bl_int_66_61 bl_int_65_61 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c62
+ bl_int_66_62 bl_int_65_62 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c63
+ bl_int_66_63 bl_int_65_63 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c64
+ bl_int_66_64 bl_int_65_64 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c65
+ bl_int_66_65 bl_int_65_65 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c66
+ bl_int_66_66 bl_int_65_66 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c67
+ bl_int_66_67 bl_int_65_67 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c68
+ bl_int_66_68 bl_int_65_68 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c69
+ bl_int_66_69 bl_int_65_69 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c70
+ bl_int_66_70 bl_int_65_70 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c71
+ bl_int_66_71 bl_int_65_71 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c72
+ bl_int_66_72 bl_int_65_72 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c73
+ bl_int_66_73 bl_int_65_73 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c74
+ bl_int_66_74 bl_int_65_74 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c75
+ bl_int_66_75 bl_int_65_75 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c76
+ bl_int_66_76 bl_int_65_76 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c77
+ bl_int_66_77 bl_int_65_77 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c78
+ bl_int_66_78 bl_int_65_78 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c79
+ bl_int_66_79 bl_int_65_79 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c80
+ bl_int_66_80 bl_int_65_80 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c81
+ bl_int_66_81 bl_int_65_81 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c82
+ bl_int_66_82 bl_int_65_82 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c83
+ bl_int_66_83 bl_int_65_83 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c84
+ bl_int_66_84 bl_int_65_84 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c85
+ bl_int_66_85 bl_int_65_85 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c86
+ bl_int_66_86 bl_int_65_86 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c87
+ bl_int_66_87 bl_int_65_87 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c88
+ bl_int_66_88 bl_int_65_88 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c89
+ bl_int_66_89 bl_int_65_89 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c90
+ bl_int_66_90 bl_int_65_90 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c91
+ bl_int_66_91 bl_int_65_91 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c92
+ bl_int_66_92 bl_int_65_92 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c93
+ bl_int_66_93 bl_int_65_93 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c94
+ bl_int_66_94 bl_int_65_94 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c95
+ bl_int_66_95 bl_int_65_95 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c96
+ bl_int_66_96 bl_int_65_96 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c97
+ bl_int_66_97 bl_int_65_97 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c98
+ bl_int_66_98 bl_int_65_98 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c99
+ bl_int_66_99 bl_int_65_99 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c100
+ bl_int_66_100 bl_int_65_100 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c101
+ bl_int_66_101 bl_int_65_101 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c102
+ bl_int_66_102 bl_int_65_102 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c103
+ bl_int_66_103 bl_int_65_103 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c104
+ bl_int_66_104 bl_int_65_104 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c105
+ bl_int_66_105 bl_int_65_105 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c106
+ bl_int_66_106 bl_int_65_106 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c107
+ bl_int_66_107 bl_int_65_107 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c108
+ bl_int_66_108 bl_int_65_108 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c109
+ bl_int_66_109 bl_int_65_109 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c110
+ bl_int_66_110 bl_int_65_110 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c111
+ bl_int_66_111 bl_int_65_111 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c112
+ bl_int_66_112 bl_int_65_112 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c113
+ bl_int_66_113 bl_int_65_113 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c114
+ bl_int_66_114 bl_int_65_114 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c115
+ bl_int_66_115 bl_int_65_115 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c116
+ bl_int_66_116 bl_int_65_116 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c117
+ bl_int_66_117 bl_int_65_117 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c118
+ bl_int_66_118 bl_int_65_118 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c119
+ bl_int_66_119 bl_int_65_119 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c120
+ bl_int_66_120 bl_int_65_120 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c121
+ bl_int_66_121 bl_int_65_121 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c122
+ bl_int_66_122 bl_int_65_122 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c123
+ bl_int_66_123 bl_int_65_123 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c124
+ bl_int_66_124 bl_int_65_124 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c125
+ bl_int_66_125 bl_int_65_125 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c126
+ bl_int_66_126 bl_int_65_126 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c127
+ bl_int_66_127 bl_int_65_127 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c128
+ bl_int_66_128 bl_int_65_128 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c129
+ bl_int_66_129 bl_int_65_129 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c130
+ bl_int_66_130 bl_int_65_130 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c131
+ bl_int_66_131 bl_int_65_131 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c132
+ bl_int_66_132 bl_int_65_132 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c133
+ bl_int_66_133 bl_int_65_133 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c134
+ bl_int_66_134 bl_int_65_134 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c135
+ bl_int_66_135 bl_int_65_135 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c136
+ bl_int_66_136 bl_int_65_136 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c137
+ bl_int_66_137 bl_int_65_137 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c138
+ bl_int_66_138 bl_int_65_138 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c139
+ bl_int_66_139 bl_int_65_139 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c140
+ bl_int_66_140 bl_int_65_140 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c141
+ bl_int_66_141 bl_int_65_141 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c142
+ bl_int_66_142 bl_int_65_142 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c143
+ bl_int_66_143 bl_int_65_143 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c144
+ bl_int_66_144 bl_int_65_144 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c145
+ bl_int_66_145 bl_int_65_145 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c146
+ bl_int_66_146 bl_int_65_146 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c147
+ bl_int_66_147 bl_int_65_147 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c148
+ bl_int_66_148 bl_int_65_148 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c149
+ bl_int_66_149 bl_int_65_149 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c150
+ bl_int_66_150 bl_int_65_150 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c151
+ bl_int_66_151 bl_int_65_151 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c152
+ bl_int_66_152 bl_int_65_152 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c153
+ bl_int_66_153 bl_int_65_153 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c154
+ bl_int_66_154 bl_int_65_154 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c155
+ bl_int_66_155 bl_int_65_155 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c156
+ bl_int_66_156 bl_int_65_156 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c157
+ bl_int_66_157 bl_int_65_157 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c158
+ bl_int_66_158 bl_int_65_158 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c159
+ bl_int_66_159 bl_int_65_159 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c160
+ bl_int_66_160 bl_int_65_160 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c161
+ bl_int_66_161 bl_int_65_161 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c162
+ bl_int_66_162 bl_int_65_162 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c163
+ bl_int_66_163 bl_int_65_163 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c164
+ bl_int_66_164 bl_int_65_164 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c165
+ bl_int_66_165 bl_int_65_165 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c166
+ bl_int_66_166 bl_int_65_166 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c167
+ bl_int_66_167 bl_int_65_167 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c168
+ bl_int_66_168 bl_int_65_168 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c169
+ bl_int_66_169 bl_int_65_169 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c170
+ bl_int_66_170 bl_int_65_170 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c171
+ bl_int_66_171 bl_int_65_171 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c172
+ bl_int_66_172 bl_int_65_172 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c173
+ bl_int_66_173 bl_int_65_173 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c174
+ bl_int_66_174 bl_int_65_174 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c175
+ bl_int_66_175 bl_int_65_175 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c176
+ bl_int_66_176 bl_int_65_176 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c177
+ bl_int_66_177 bl_int_65_177 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c178
+ bl_int_66_178 bl_int_65_178 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c179
+ bl_int_66_179 bl_int_65_179 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c180
+ bl_int_66_180 bl_int_65_180 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c181
+ bl_int_66_181 bl_int_65_181 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c182
+ bl_int_66_182 bl_int_65_182 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r66_c183
+ bl_int_66_183 bl_int_65_183 wl_0_66 gnd
+ sram_rom_base_one_cell
Xbit_r67_c0
+ bl_int_67_0 bl_int_66_0 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c1
+ bl_int_67_1 bl_int_66_1 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c2
+ bl_int_67_2 bl_int_66_2 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c3
+ bl_int_67_3 bl_int_66_3 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c4
+ bl_int_67_4 bl_int_66_4 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c5
+ bl_int_67_5 bl_int_66_5 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c6
+ bl_int_67_6 bl_int_66_6 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c7
+ bl_int_67_7 bl_int_66_7 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c8
+ bl_int_67_8 bl_int_66_8 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c9
+ bl_int_67_9 bl_int_66_9 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c10
+ bl_int_67_10 bl_int_66_10 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c11
+ bl_int_67_11 bl_int_66_11 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c12
+ bl_int_67_12 bl_int_66_12 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c13
+ bl_int_67_13 bl_int_66_13 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c14
+ bl_int_67_14 bl_int_66_14 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c15
+ bl_int_67_15 bl_int_66_15 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c16
+ bl_int_67_16 bl_int_66_16 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c17
+ bl_int_67_17 bl_int_66_17 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c18
+ bl_int_67_18 bl_int_66_18 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c19
+ bl_int_67_19 bl_int_66_19 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c20
+ bl_int_67_20 bl_int_66_20 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c21
+ bl_int_67_21 bl_int_66_21 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c22
+ bl_int_67_22 bl_int_66_22 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c23
+ bl_int_67_23 bl_int_66_23 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c24
+ bl_int_67_24 bl_int_66_24 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c25
+ bl_int_67_25 bl_int_66_25 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c26
+ bl_int_67_26 bl_int_66_26 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c27
+ bl_int_67_27 bl_int_66_27 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c28
+ bl_int_67_28 bl_int_66_28 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c29
+ bl_int_67_29 bl_int_66_29 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c30
+ bl_int_67_30 bl_int_66_30 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c31
+ bl_int_67_31 bl_int_66_31 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c32
+ bl_int_67_32 bl_int_66_32 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c33
+ bl_int_67_33 bl_int_66_33 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c34
+ bl_int_67_34 bl_int_66_34 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c35
+ bl_int_67_35 bl_int_66_35 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c36
+ bl_int_67_36 bl_int_66_36 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c37
+ bl_int_67_37 bl_int_66_37 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c38
+ bl_int_67_38 bl_int_66_38 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c39
+ bl_int_67_39 bl_int_66_39 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c40
+ bl_int_67_40 bl_int_66_40 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c41
+ bl_int_67_41 bl_int_66_41 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c42
+ bl_int_67_42 bl_int_66_42 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c43
+ bl_int_67_43 bl_int_66_43 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c44
+ bl_int_67_44 bl_int_66_44 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c45
+ bl_int_67_45 bl_int_66_45 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c46
+ bl_int_67_46 bl_int_66_46 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c47
+ bl_int_67_47 bl_int_66_47 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c48
+ bl_int_67_48 bl_int_66_48 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c49
+ bl_int_67_49 bl_int_66_49 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c50
+ bl_int_67_50 bl_int_66_50 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c51
+ bl_int_67_51 bl_int_66_51 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c52
+ bl_int_67_52 bl_int_66_52 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c53
+ bl_int_67_53 bl_int_66_53 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c54
+ bl_int_67_54 bl_int_66_54 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c55
+ bl_int_67_55 bl_int_66_55 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c56
+ bl_int_67_56 bl_int_66_56 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c57
+ bl_int_67_57 bl_int_66_57 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c58
+ bl_int_67_58 bl_int_66_58 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c59
+ bl_int_67_59 bl_int_66_59 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c60
+ bl_int_67_60 bl_int_66_60 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c61
+ bl_int_67_61 bl_int_66_61 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c62
+ bl_int_67_62 bl_int_66_62 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c63
+ bl_int_67_63 bl_int_66_63 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c64
+ bl_int_67_64 bl_int_66_64 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c65
+ bl_int_67_65 bl_int_66_65 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c66
+ bl_int_67_66 bl_int_66_66 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c67
+ bl_int_67_67 bl_int_66_67 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c68
+ bl_int_67_68 bl_int_66_68 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c69
+ bl_int_67_69 bl_int_66_69 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c70
+ bl_int_67_70 bl_int_66_70 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c71
+ bl_int_67_71 bl_int_66_71 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c72
+ bl_int_67_72 bl_int_66_72 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c73
+ bl_int_67_73 bl_int_66_73 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c74
+ bl_int_67_74 bl_int_66_74 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c75
+ bl_int_67_75 bl_int_66_75 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c76
+ bl_int_67_76 bl_int_66_76 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c77
+ bl_int_67_77 bl_int_66_77 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c78
+ bl_int_67_78 bl_int_66_78 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c79
+ bl_int_67_79 bl_int_66_79 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c80
+ bl_int_67_80 bl_int_66_80 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c81
+ bl_int_67_81 bl_int_66_81 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c82
+ bl_int_67_82 bl_int_66_82 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c83
+ bl_int_67_83 bl_int_66_83 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c84
+ bl_int_67_84 bl_int_66_84 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c85
+ bl_int_67_85 bl_int_66_85 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c86
+ bl_int_67_86 bl_int_66_86 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c87
+ bl_int_67_87 bl_int_66_87 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c88
+ bl_int_67_88 bl_int_66_88 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c89
+ bl_int_67_89 bl_int_66_89 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c90
+ bl_int_67_90 bl_int_66_90 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c91
+ bl_int_67_91 bl_int_66_91 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c92
+ bl_int_67_92 bl_int_66_92 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c93
+ bl_int_67_93 bl_int_66_93 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c94
+ bl_int_67_94 bl_int_66_94 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c95
+ bl_int_67_95 bl_int_66_95 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c96
+ bl_int_67_96 bl_int_66_96 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c97
+ bl_int_67_97 bl_int_66_97 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c98
+ bl_int_67_98 bl_int_66_98 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c99
+ bl_int_67_99 bl_int_66_99 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c100
+ bl_int_67_100 bl_int_66_100 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c101
+ bl_int_67_101 bl_int_66_101 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c102
+ bl_int_67_102 bl_int_66_102 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c103
+ bl_int_67_103 bl_int_66_103 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c104
+ bl_int_67_104 bl_int_66_104 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c105
+ bl_int_67_105 bl_int_66_105 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c106
+ bl_int_67_106 bl_int_66_106 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c107
+ bl_int_67_107 bl_int_66_107 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c108
+ bl_int_67_108 bl_int_66_108 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c109
+ bl_int_67_109 bl_int_66_109 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c110
+ bl_int_67_110 bl_int_66_110 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c111
+ bl_int_67_111 bl_int_66_111 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c112
+ bl_int_67_112 bl_int_66_112 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c113
+ bl_int_67_113 bl_int_66_113 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c114
+ bl_int_67_114 bl_int_66_114 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c115
+ bl_int_67_115 bl_int_66_115 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c116
+ bl_int_67_116 bl_int_66_116 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c117
+ bl_int_67_117 bl_int_66_117 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c118
+ bl_int_67_118 bl_int_66_118 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c119
+ bl_int_67_119 bl_int_66_119 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c120
+ bl_int_67_120 bl_int_66_120 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c121
+ bl_int_67_121 bl_int_66_121 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c122
+ bl_int_67_122 bl_int_66_122 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c123
+ bl_int_67_123 bl_int_66_123 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c124
+ bl_int_67_124 bl_int_66_124 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c125
+ bl_int_67_125 bl_int_66_125 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c126
+ bl_int_67_126 bl_int_66_126 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c127
+ bl_int_67_127 bl_int_66_127 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c128
+ bl_int_67_128 bl_int_66_128 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c129
+ bl_int_67_129 bl_int_66_129 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c130
+ bl_int_67_130 bl_int_66_130 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c131
+ bl_int_67_131 bl_int_66_131 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c132
+ bl_int_67_132 bl_int_66_132 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c133
+ bl_int_67_133 bl_int_66_133 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c134
+ bl_int_67_134 bl_int_66_134 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c135
+ bl_int_67_135 bl_int_66_135 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c136
+ bl_int_67_136 bl_int_66_136 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c137
+ bl_int_67_137 bl_int_66_137 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c138
+ bl_int_67_138 bl_int_66_138 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c139
+ bl_int_67_139 bl_int_66_139 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c140
+ bl_int_67_140 bl_int_66_140 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c141
+ bl_int_67_141 bl_int_66_141 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c142
+ bl_int_67_142 bl_int_66_142 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c143
+ bl_int_67_143 bl_int_66_143 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c144
+ bl_int_67_144 bl_int_66_144 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c145
+ bl_int_67_145 bl_int_66_145 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c146
+ bl_int_67_146 bl_int_66_146 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c147
+ bl_int_67_147 bl_int_66_147 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c148
+ bl_int_67_148 bl_int_66_148 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c149
+ bl_int_67_149 bl_int_66_149 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c150
+ bl_int_67_150 bl_int_66_150 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c151
+ bl_int_67_151 bl_int_66_151 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c152
+ bl_int_67_152 bl_int_66_152 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c153
+ bl_int_67_153 bl_int_66_153 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c154
+ bl_int_67_154 bl_int_66_154 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c155
+ bl_int_67_155 bl_int_66_155 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c156
+ bl_int_67_156 bl_int_66_156 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c157
+ bl_int_67_157 bl_int_66_157 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c158
+ bl_int_67_158 bl_int_66_158 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c159
+ bl_int_67_159 bl_int_66_159 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c160
+ bl_int_67_160 bl_int_66_160 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c161
+ bl_int_67_161 bl_int_66_161 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c162
+ bl_int_67_162 bl_int_66_162 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c163
+ bl_int_67_163 bl_int_66_163 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c164
+ bl_int_67_164 bl_int_66_164 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c165
+ bl_int_67_165 bl_int_66_165 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c166
+ bl_int_67_166 bl_int_66_166 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c167
+ bl_int_67_167 bl_int_66_167 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c168
+ bl_int_67_168 bl_int_66_168 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c169
+ bl_int_67_169 bl_int_66_169 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c170
+ bl_int_67_170 bl_int_66_170 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c171
+ bl_int_67_171 bl_int_66_171 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c172
+ bl_int_67_172 bl_int_66_172 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c173
+ bl_int_67_173 bl_int_66_173 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c174
+ bl_int_67_174 bl_int_66_174 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c175
+ bl_int_67_175 bl_int_66_175 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c176
+ bl_int_67_176 bl_int_66_176 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c177
+ bl_int_67_177 bl_int_66_177 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c178
+ bl_int_67_178 bl_int_66_178 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c179
+ bl_int_67_179 bl_int_66_179 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c180
+ bl_int_67_180 bl_int_66_180 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c181
+ bl_int_67_181 bl_int_66_181 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c182
+ bl_int_67_182 bl_int_66_182 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r67_c183
+ bl_int_67_183 bl_int_66_183 wl_0_67 gnd
+ sram_rom_base_one_cell
Xbit_r68_c0
+ bl_int_68_0 bl_int_67_0 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c1
+ bl_int_68_1 bl_int_67_1 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c2
+ bl_int_68_2 bl_int_67_2 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c3
+ bl_int_68_3 bl_int_67_3 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c4
+ bl_int_68_4 bl_int_67_4 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c5
+ bl_int_68_5 bl_int_67_5 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c6
+ bl_int_68_6 bl_int_67_6 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c7
+ bl_int_68_7 bl_int_67_7 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c8
+ bl_int_68_8 bl_int_67_8 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c9
+ bl_int_68_9 bl_int_67_9 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c10
+ bl_int_68_10 bl_int_67_10 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c11
+ bl_int_68_11 bl_int_67_11 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c12
+ bl_int_68_12 bl_int_67_12 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c13
+ bl_int_68_13 bl_int_67_13 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c14
+ bl_int_68_14 bl_int_67_14 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c15
+ bl_int_68_15 bl_int_67_15 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c16
+ bl_int_68_16 bl_int_67_16 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c17
+ bl_int_68_17 bl_int_67_17 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c18
+ bl_int_68_18 bl_int_67_18 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c19
+ bl_int_68_19 bl_int_67_19 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c20
+ bl_int_68_20 bl_int_67_20 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c21
+ bl_int_68_21 bl_int_67_21 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c22
+ bl_int_68_22 bl_int_67_22 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c23
+ bl_int_68_23 bl_int_67_23 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c24
+ bl_int_68_24 bl_int_67_24 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c25
+ bl_int_68_25 bl_int_67_25 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c26
+ bl_int_68_26 bl_int_67_26 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c27
+ bl_int_68_27 bl_int_67_27 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c28
+ bl_int_68_28 bl_int_67_28 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c29
+ bl_int_68_29 bl_int_67_29 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c30
+ bl_int_68_30 bl_int_67_30 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c31
+ bl_int_68_31 bl_int_67_31 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c32
+ bl_int_68_32 bl_int_67_32 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c33
+ bl_int_68_33 bl_int_67_33 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c34
+ bl_int_68_34 bl_int_67_34 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c35
+ bl_int_68_35 bl_int_67_35 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c36
+ bl_int_68_36 bl_int_67_36 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c37
+ bl_int_68_37 bl_int_67_37 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c38
+ bl_int_68_38 bl_int_67_38 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c39
+ bl_int_68_39 bl_int_67_39 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c40
+ bl_int_68_40 bl_int_67_40 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c41
+ bl_int_68_41 bl_int_67_41 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c42
+ bl_int_68_42 bl_int_67_42 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c43
+ bl_int_68_43 bl_int_67_43 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c44
+ bl_int_68_44 bl_int_67_44 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c45
+ bl_int_68_45 bl_int_67_45 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c46
+ bl_int_68_46 bl_int_67_46 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c47
+ bl_int_68_47 bl_int_67_47 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c48
+ bl_int_68_48 bl_int_67_48 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c49
+ bl_int_68_49 bl_int_67_49 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c50
+ bl_int_68_50 bl_int_67_50 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c51
+ bl_int_68_51 bl_int_67_51 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c52
+ bl_int_68_52 bl_int_67_52 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c53
+ bl_int_68_53 bl_int_67_53 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c54
+ bl_int_68_54 bl_int_67_54 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c55
+ bl_int_68_55 bl_int_67_55 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c56
+ bl_int_68_56 bl_int_67_56 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c57
+ bl_int_68_57 bl_int_67_57 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c58
+ bl_int_68_58 bl_int_67_58 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c59
+ bl_int_68_59 bl_int_67_59 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c60
+ bl_int_68_60 bl_int_67_60 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c61
+ bl_int_68_61 bl_int_67_61 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c62
+ bl_int_68_62 bl_int_67_62 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c63
+ bl_int_68_63 bl_int_67_63 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c64
+ bl_int_68_64 bl_int_67_64 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c65
+ bl_int_68_65 bl_int_67_65 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c66
+ bl_int_68_66 bl_int_67_66 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c67
+ bl_int_68_67 bl_int_67_67 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c68
+ bl_int_68_68 bl_int_67_68 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c69
+ bl_int_68_69 bl_int_67_69 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c70
+ bl_int_68_70 bl_int_67_70 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c71
+ bl_int_68_71 bl_int_67_71 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c72
+ bl_int_68_72 bl_int_67_72 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c73
+ bl_int_68_73 bl_int_67_73 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c74
+ bl_int_68_74 bl_int_67_74 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c75
+ bl_int_68_75 bl_int_67_75 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c76
+ bl_int_68_76 bl_int_67_76 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c77
+ bl_int_68_77 bl_int_67_77 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c78
+ bl_int_68_78 bl_int_67_78 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c79
+ bl_int_68_79 bl_int_67_79 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c80
+ bl_int_68_80 bl_int_67_80 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c81
+ bl_int_68_81 bl_int_67_81 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c82
+ bl_int_68_82 bl_int_67_82 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c83
+ bl_int_68_83 bl_int_67_83 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c84
+ bl_int_68_84 bl_int_67_84 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c85
+ bl_int_68_85 bl_int_67_85 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c86
+ bl_int_68_86 bl_int_67_86 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c87
+ bl_int_68_87 bl_int_67_87 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c88
+ bl_int_68_88 bl_int_67_88 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c89
+ bl_int_68_89 bl_int_67_89 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c90
+ bl_int_68_90 bl_int_67_90 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c91
+ bl_int_68_91 bl_int_67_91 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c92
+ bl_int_68_92 bl_int_67_92 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c93
+ bl_int_68_93 bl_int_67_93 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c94
+ bl_int_68_94 bl_int_67_94 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c95
+ bl_int_68_95 bl_int_67_95 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c96
+ bl_int_68_96 bl_int_67_96 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c97
+ bl_int_68_97 bl_int_67_97 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c98
+ bl_int_68_98 bl_int_67_98 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c99
+ bl_int_68_99 bl_int_67_99 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c100
+ bl_int_68_100 bl_int_67_100 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c101
+ bl_int_68_101 bl_int_67_101 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c102
+ bl_int_68_102 bl_int_67_102 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c103
+ bl_int_68_103 bl_int_67_103 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c104
+ bl_int_68_104 bl_int_67_104 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c105
+ bl_int_68_105 bl_int_67_105 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c106
+ bl_int_68_106 bl_int_67_106 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c107
+ bl_int_68_107 bl_int_67_107 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c108
+ bl_int_68_108 bl_int_67_108 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c109
+ bl_int_68_109 bl_int_67_109 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c110
+ bl_int_68_110 bl_int_67_110 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c111
+ bl_int_68_111 bl_int_67_111 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c112
+ bl_int_68_112 bl_int_67_112 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c113
+ bl_int_68_113 bl_int_67_113 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c114
+ bl_int_68_114 bl_int_67_114 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c115
+ bl_int_68_115 bl_int_67_115 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c116
+ bl_int_68_116 bl_int_67_116 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c117
+ bl_int_68_117 bl_int_67_117 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c118
+ bl_int_68_118 bl_int_67_118 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c119
+ bl_int_68_119 bl_int_67_119 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c120
+ bl_int_68_120 bl_int_67_120 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c121
+ bl_int_68_121 bl_int_67_121 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c122
+ bl_int_68_122 bl_int_67_122 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c123
+ bl_int_68_123 bl_int_67_123 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c124
+ bl_int_68_124 bl_int_67_124 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c125
+ bl_int_68_125 bl_int_67_125 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c126
+ bl_int_68_126 bl_int_67_126 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c127
+ bl_int_68_127 bl_int_67_127 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c128
+ bl_int_68_128 bl_int_67_128 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c129
+ bl_int_68_129 bl_int_67_129 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c130
+ bl_int_68_130 bl_int_67_130 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c131
+ bl_int_68_131 bl_int_67_131 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c132
+ bl_int_68_132 bl_int_67_132 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c133
+ bl_int_68_133 bl_int_67_133 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c134
+ bl_int_68_134 bl_int_67_134 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c135
+ bl_int_68_135 bl_int_67_135 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c136
+ bl_int_68_136 bl_int_67_136 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c137
+ bl_int_68_137 bl_int_67_137 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c138
+ bl_int_68_138 bl_int_67_138 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c139
+ bl_int_68_139 bl_int_67_139 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c140
+ bl_int_68_140 bl_int_67_140 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c141
+ bl_int_68_141 bl_int_67_141 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c142
+ bl_int_68_142 bl_int_67_142 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c143
+ bl_int_68_143 bl_int_67_143 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c144
+ bl_int_68_144 bl_int_67_144 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c145
+ bl_int_68_145 bl_int_67_145 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c146
+ bl_int_68_146 bl_int_67_146 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c147
+ bl_int_68_147 bl_int_67_147 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c148
+ bl_int_68_148 bl_int_67_148 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c149
+ bl_int_68_149 bl_int_67_149 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c150
+ bl_int_68_150 bl_int_67_150 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c151
+ bl_int_68_151 bl_int_67_151 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c152
+ bl_int_68_152 bl_int_67_152 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c153
+ bl_int_68_153 bl_int_67_153 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c154
+ bl_int_68_154 bl_int_67_154 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c155
+ bl_int_68_155 bl_int_67_155 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c156
+ bl_int_68_156 bl_int_67_156 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c157
+ bl_int_68_157 bl_int_67_157 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c158
+ bl_int_68_158 bl_int_67_158 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c159
+ bl_int_68_159 bl_int_67_159 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c160
+ bl_int_68_160 bl_int_67_160 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c161
+ bl_int_68_161 bl_int_67_161 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c162
+ bl_int_68_162 bl_int_67_162 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c163
+ bl_int_68_163 bl_int_67_163 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c164
+ bl_int_68_164 bl_int_67_164 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c165
+ bl_int_68_165 bl_int_67_165 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c166
+ bl_int_68_166 bl_int_67_166 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c167
+ bl_int_68_167 bl_int_67_167 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c168
+ bl_int_68_168 bl_int_67_168 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c169
+ bl_int_68_169 bl_int_67_169 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c170
+ bl_int_68_170 bl_int_67_170 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c171
+ bl_int_68_171 bl_int_67_171 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c172
+ bl_int_68_172 bl_int_67_172 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c173
+ bl_int_68_173 bl_int_67_173 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c174
+ bl_int_68_174 bl_int_67_174 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c175
+ bl_int_68_175 bl_int_67_175 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c176
+ bl_int_68_176 bl_int_67_176 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c177
+ bl_int_68_177 bl_int_67_177 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c178
+ bl_int_68_178 bl_int_67_178 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c179
+ bl_int_68_179 bl_int_67_179 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c180
+ bl_int_68_180 bl_int_67_180 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c181
+ bl_int_68_181 bl_int_67_181 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c182
+ bl_int_68_182 bl_int_67_182 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r68_c183
+ bl_int_68_183 bl_int_67_183 wl_0_68 gnd
+ sram_rom_base_one_cell
Xbit_r69_c0
+ bl_int_69_0 bl_int_68_0 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c1
+ bl_int_69_1 bl_int_68_1 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c2
+ bl_int_69_2 bl_int_68_2 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c3
+ bl_int_69_3 bl_int_68_3 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c4
+ bl_int_69_4 bl_int_68_4 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c5
+ bl_int_69_5 bl_int_68_5 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c6
+ bl_int_69_6 bl_int_68_6 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c7
+ bl_int_69_7 bl_int_68_7 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c8
+ bl_int_69_8 bl_int_68_8 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c9
+ bl_int_69_9 bl_int_68_9 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c10
+ bl_int_69_10 bl_int_68_10 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c11
+ bl_int_69_11 bl_int_68_11 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c12
+ bl_int_69_12 bl_int_68_12 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c13
+ bl_int_69_13 bl_int_68_13 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c14
+ bl_int_69_14 bl_int_68_14 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c15
+ bl_int_69_15 bl_int_68_15 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c16
+ bl_int_69_16 bl_int_68_16 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c17
+ bl_int_69_17 bl_int_68_17 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c18
+ bl_int_69_18 bl_int_68_18 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c19
+ bl_int_69_19 bl_int_68_19 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c20
+ bl_int_69_20 bl_int_68_20 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c21
+ bl_int_69_21 bl_int_68_21 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c22
+ bl_int_69_22 bl_int_68_22 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c23
+ bl_int_69_23 bl_int_68_23 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c24
+ bl_int_69_24 bl_int_68_24 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c25
+ bl_int_69_25 bl_int_68_25 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c26
+ bl_int_69_26 bl_int_68_26 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c27
+ bl_int_69_27 bl_int_68_27 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c28
+ bl_int_69_28 bl_int_68_28 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c29
+ bl_int_69_29 bl_int_68_29 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c30
+ bl_int_69_30 bl_int_68_30 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c31
+ bl_int_69_31 bl_int_68_31 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c32
+ bl_int_69_32 bl_int_68_32 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c33
+ bl_int_69_33 bl_int_68_33 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c34
+ bl_int_69_34 bl_int_68_34 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c35
+ bl_int_69_35 bl_int_68_35 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c36
+ bl_int_69_36 bl_int_68_36 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c37
+ bl_int_69_37 bl_int_68_37 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c38
+ bl_int_69_38 bl_int_68_38 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c39
+ bl_int_69_39 bl_int_68_39 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c40
+ bl_int_69_40 bl_int_68_40 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c41
+ bl_int_69_41 bl_int_68_41 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c42
+ bl_int_69_42 bl_int_68_42 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c43
+ bl_int_69_43 bl_int_68_43 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c44
+ bl_int_69_44 bl_int_68_44 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c45
+ bl_int_69_45 bl_int_68_45 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c46
+ bl_int_69_46 bl_int_68_46 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c47
+ bl_int_69_47 bl_int_68_47 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c48
+ bl_int_69_48 bl_int_68_48 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c49
+ bl_int_69_49 bl_int_68_49 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c50
+ bl_int_69_50 bl_int_68_50 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c51
+ bl_int_69_51 bl_int_68_51 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c52
+ bl_int_69_52 bl_int_68_52 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c53
+ bl_int_69_53 bl_int_68_53 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c54
+ bl_int_69_54 bl_int_68_54 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c55
+ bl_int_69_55 bl_int_68_55 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c56
+ bl_int_69_56 bl_int_68_56 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c57
+ bl_int_69_57 bl_int_68_57 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c58
+ bl_int_69_58 bl_int_68_58 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c59
+ bl_int_69_59 bl_int_68_59 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c60
+ bl_int_69_60 bl_int_68_60 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c61
+ bl_int_69_61 bl_int_68_61 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c62
+ bl_int_69_62 bl_int_68_62 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c63
+ bl_int_69_63 bl_int_68_63 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c64
+ bl_int_69_64 bl_int_68_64 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c65
+ bl_int_69_65 bl_int_68_65 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c66
+ bl_int_69_66 bl_int_68_66 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c67
+ bl_int_69_67 bl_int_68_67 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c68
+ bl_int_69_68 bl_int_68_68 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c69
+ bl_int_69_69 bl_int_68_69 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c70
+ bl_int_69_70 bl_int_68_70 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c71
+ bl_int_69_71 bl_int_68_71 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c72
+ bl_int_69_72 bl_int_68_72 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c73
+ bl_int_69_73 bl_int_68_73 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c74
+ bl_int_69_74 bl_int_68_74 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c75
+ bl_int_69_75 bl_int_68_75 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c76
+ bl_int_69_76 bl_int_68_76 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c77
+ bl_int_69_77 bl_int_68_77 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c78
+ bl_int_69_78 bl_int_68_78 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c79
+ bl_int_69_79 bl_int_68_79 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c80
+ bl_int_69_80 bl_int_68_80 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c81
+ bl_int_69_81 bl_int_68_81 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c82
+ bl_int_69_82 bl_int_68_82 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c83
+ bl_int_69_83 bl_int_68_83 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c84
+ bl_int_69_84 bl_int_68_84 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c85
+ bl_int_69_85 bl_int_68_85 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c86
+ bl_int_69_86 bl_int_68_86 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c87
+ bl_int_69_87 bl_int_68_87 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c88
+ bl_int_69_88 bl_int_68_88 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c89
+ bl_int_69_89 bl_int_68_89 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c90
+ bl_int_69_90 bl_int_68_90 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c91
+ bl_int_69_91 bl_int_68_91 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c92
+ bl_int_69_92 bl_int_68_92 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c93
+ bl_int_69_93 bl_int_68_93 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c94
+ bl_int_69_94 bl_int_68_94 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c95
+ bl_int_69_95 bl_int_68_95 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c96
+ bl_int_69_96 bl_int_68_96 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c97
+ bl_int_69_97 bl_int_68_97 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c98
+ bl_int_69_98 bl_int_68_98 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c99
+ bl_int_69_99 bl_int_68_99 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c100
+ bl_int_69_100 bl_int_68_100 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c101
+ bl_int_69_101 bl_int_68_101 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c102
+ bl_int_69_102 bl_int_68_102 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c103
+ bl_int_69_103 bl_int_68_103 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c104
+ bl_int_69_104 bl_int_68_104 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c105
+ bl_int_69_105 bl_int_68_105 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c106
+ bl_int_69_106 bl_int_68_106 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c107
+ bl_int_69_107 bl_int_68_107 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c108
+ bl_int_69_108 bl_int_68_108 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c109
+ bl_int_69_109 bl_int_68_109 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c110
+ bl_int_69_110 bl_int_68_110 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c111
+ bl_int_69_111 bl_int_68_111 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c112
+ bl_int_69_112 bl_int_68_112 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c113
+ bl_int_69_113 bl_int_68_113 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c114
+ bl_int_69_114 bl_int_68_114 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c115
+ bl_int_69_115 bl_int_68_115 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c116
+ bl_int_69_116 bl_int_68_116 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c117
+ bl_int_69_117 bl_int_68_117 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c118
+ bl_int_69_118 bl_int_68_118 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c119
+ bl_int_69_119 bl_int_68_119 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c120
+ bl_int_69_120 bl_int_68_120 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c121
+ bl_int_69_121 bl_int_68_121 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c122
+ bl_int_69_122 bl_int_68_122 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c123
+ bl_int_69_123 bl_int_68_123 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c124
+ bl_int_69_124 bl_int_68_124 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c125
+ bl_int_69_125 bl_int_68_125 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c126
+ bl_int_69_126 bl_int_68_126 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c127
+ bl_int_69_127 bl_int_68_127 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c128
+ bl_int_69_128 bl_int_68_128 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c129
+ bl_int_69_129 bl_int_68_129 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c130
+ bl_int_69_130 bl_int_68_130 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c131
+ bl_int_69_131 bl_int_68_131 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c132
+ bl_int_69_132 bl_int_68_132 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c133
+ bl_int_69_133 bl_int_68_133 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c134
+ bl_int_69_134 bl_int_68_134 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c135
+ bl_int_69_135 bl_int_68_135 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c136
+ bl_int_69_136 bl_int_68_136 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c137
+ bl_int_69_137 bl_int_68_137 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c138
+ bl_int_69_138 bl_int_68_138 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c139
+ bl_int_69_139 bl_int_68_139 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c140
+ bl_int_69_140 bl_int_68_140 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c141
+ bl_int_69_141 bl_int_68_141 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c142
+ bl_int_69_142 bl_int_68_142 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c143
+ bl_int_69_143 bl_int_68_143 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c144
+ bl_int_69_144 bl_int_68_144 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c145
+ bl_int_69_145 bl_int_68_145 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c146
+ bl_int_69_146 bl_int_68_146 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c147
+ bl_int_69_147 bl_int_68_147 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c148
+ bl_int_69_148 bl_int_68_148 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c149
+ bl_int_69_149 bl_int_68_149 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c150
+ bl_int_69_150 bl_int_68_150 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c151
+ bl_int_69_151 bl_int_68_151 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c152
+ bl_int_69_152 bl_int_68_152 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c153
+ bl_int_69_153 bl_int_68_153 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c154
+ bl_int_69_154 bl_int_68_154 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c155
+ bl_int_69_155 bl_int_68_155 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c156
+ bl_int_69_156 bl_int_68_156 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c157
+ bl_int_69_157 bl_int_68_157 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c158
+ bl_int_69_158 bl_int_68_158 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c159
+ bl_int_69_159 bl_int_68_159 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c160
+ bl_int_69_160 bl_int_68_160 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c161
+ bl_int_69_161 bl_int_68_161 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c162
+ bl_int_69_162 bl_int_68_162 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c163
+ bl_int_69_163 bl_int_68_163 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c164
+ bl_int_69_164 bl_int_68_164 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c165
+ bl_int_69_165 bl_int_68_165 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c166
+ bl_int_69_166 bl_int_68_166 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c167
+ bl_int_69_167 bl_int_68_167 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c168
+ bl_int_69_168 bl_int_68_168 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c169
+ bl_int_69_169 bl_int_68_169 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c170
+ bl_int_69_170 bl_int_68_170 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c171
+ bl_int_69_171 bl_int_68_171 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c172
+ bl_int_69_172 bl_int_68_172 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c173
+ bl_int_69_173 bl_int_68_173 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c174
+ bl_int_69_174 bl_int_68_174 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c175
+ bl_int_69_175 bl_int_68_175 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c176
+ bl_int_69_176 bl_int_68_176 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c177
+ bl_int_69_177 bl_int_68_177 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c178
+ bl_int_69_178 bl_int_68_178 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c179
+ bl_int_69_179 bl_int_68_179 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c180
+ bl_int_69_180 bl_int_68_180 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c181
+ bl_int_69_181 bl_int_68_181 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c182
+ bl_int_69_182 bl_int_68_182 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r69_c183
+ bl_int_69_183 bl_int_68_183 wl_0_69 gnd
+ sram_rom_base_one_cell
Xbit_r70_c0
+ bl_int_70_0 bl_int_69_0 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c1
+ bl_int_70_1 bl_int_69_1 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c2
+ bl_int_70_2 bl_int_69_2 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c3
+ bl_int_70_3 bl_int_69_3 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c4
+ bl_int_70_4 bl_int_69_4 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c5
+ bl_int_70_5 bl_int_69_5 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c6
+ bl_int_70_6 bl_int_69_6 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c7
+ bl_int_70_7 bl_int_69_7 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c8
+ bl_int_70_8 bl_int_69_8 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c9
+ bl_int_70_9 bl_int_69_9 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c10
+ bl_int_70_10 bl_int_69_10 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c11
+ bl_int_70_11 bl_int_69_11 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c12
+ bl_int_70_12 bl_int_69_12 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c13
+ bl_int_70_13 bl_int_69_13 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c14
+ bl_int_70_14 bl_int_69_14 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c15
+ bl_int_70_15 bl_int_69_15 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c16
+ bl_int_70_16 bl_int_69_16 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c17
+ bl_int_70_17 bl_int_69_17 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c18
+ bl_int_70_18 bl_int_69_18 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c19
+ bl_int_70_19 bl_int_69_19 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c20
+ bl_int_70_20 bl_int_69_20 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c21
+ bl_int_70_21 bl_int_69_21 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c22
+ bl_int_70_22 bl_int_69_22 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c23
+ bl_int_70_23 bl_int_69_23 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c24
+ bl_int_70_24 bl_int_69_24 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c25
+ bl_int_70_25 bl_int_69_25 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c26
+ bl_int_70_26 bl_int_69_26 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c27
+ bl_int_70_27 bl_int_69_27 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c28
+ bl_int_70_28 bl_int_69_28 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c29
+ bl_int_70_29 bl_int_69_29 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c30
+ bl_int_70_30 bl_int_69_30 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c31
+ bl_int_70_31 bl_int_69_31 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c32
+ bl_int_70_32 bl_int_69_32 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c33
+ bl_int_70_33 bl_int_69_33 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c34
+ bl_int_70_34 bl_int_69_34 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c35
+ bl_int_70_35 bl_int_69_35 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c36
+ bl_int_70_36 bl_int_69_36 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c37
+ bl_int_70_37 bl_int_69_37 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c38
+ bl_int_70_38 bl_int_69_38 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c39
+ bl_int_70_39 bl_int_69_39 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c40
+ bl_int_70_40 bl_int_69_40 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c41
+ bl_int_70_41 bl_int_69_41 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c42
+ bl_int_70_42 bl_int_69_42 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c43
+ bl_int_70_43 bl_int_69_43 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c44
+ bl_int_70_44 bl_int_69_44 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c45
+ bl_int_70_45 bl_int_69_45 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c46
+ bl_int_70_46 bl_int_69_46 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c47
+ bl_int_70_47 bl_int_69_47 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c48
+ bl_int_70_48 bl_int_69_48 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c49
+ bl_int_70_49 bl_int_69_49 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c50
+ bl_int_70_50 bl_int_69_50 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c51
+ bl_int_70_51 bl_int_69_51 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c52
+ bl_int_70_52 bl_int_69_52 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c53
+ bl_int_70_53 bl_int_69_53 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c54
+ bl_int_70_54 bl_int_69_54 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c55
+ bl_int_70_55 bl_int_69_55 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c56
+ bl_int_70_56 bl_int_69_56 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c57
+ bl_int_70_57 bl_int_69_57 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c58
+ bl_int_70_58 bl_int_69_58 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c59
+ bl_int_70_59 bl_int_69_59 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c60
+ bl_int_70_60 bl_int_69_60 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c61
+ bl_int_70_61 bl_int_69_61 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c62
+ bl_int_70_62 bl_int_69_62 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c63
+ bl_int_70_63 bl_int_69_63 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c64
+ bl_int_70_64 bl_int_69_64 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c65
+ bl_int_70_65 bl_int_69_65 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c66
+ bl_int_70_66 bl_int_69_66 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c67
+ bl_int_70_67 bl_int_69_67 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c68
+ bl_int_70_68 bl_int_69_68 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c69
+ bl_int_70_69 bl_int_69_69 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c70
+ bl_int_70_70 bl_int_69_70 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c71
+ bl_int_70_71 bl_int_69_71 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c72
+ bl_int_70_72 bl_int_69_72 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c73
+ bl_int_70_73 bl_int_69_73 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c74
+ bl_int_70_74 bl_int_69_74 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c75
+ bl_int_70_75 bl_int_69_75 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c76
+ bl_int_70_76 bl_int_69_76 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c77
+ bl_int_70_77 bl_int_69_77 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c78
+ bl_int_70_78 bl_int_69_78 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c79
+ bl_int_70_79 bl_int_69_79 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c80
+ bl_int_70_80 bl_int_69_80 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c81
+ bl_int_70_81 bl_int_69_81 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c82
+ bl_int_70_82 bl_int_69_82 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c83
+ bl_int_70_83 bl_int_69_83 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c84
+ bl_int_70_84 bl_int_69_84 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c85
+ bl_int_70_85 bl_int_69_85 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c86
+ bl_int_70_86 bl_int_69_86 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c87
+ bl_int_70_87 bl_int_69_87 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c88
+ bl_int_70_88 bl_int_69_88 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c89
+ bl_int_70_89 bl_int_69_89 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c90
+ bl_int_70_90 bl_int_69_90 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c91
+ bl_int_70_91 bl_int_69_91 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c92
+ bl_int_70_92 bl_int_69_92 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c93
+ bl_int_70_93 bl_int_69_93 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c94
+ bl_int_70_94 bl_int_69_94 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c95
+ bl_int_70_95 bl_int_69_95 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c96
+ bl_int_70_96 bl_int_69_96 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c97
+ bl_int_70_97 bl_int_69_97 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c98
+ bl_int_70_98 bl_int_69_98 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c99
+ bl_int_70_99 bl_int_69_99 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c100
+ bl_int_70_100 bl_int_69_100 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c101
+ bl_int_70_101 bl_int_69_101 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c102
+ bl_int_70_102 bl_int_69_102 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c103
+ bl_int_70_103 bl_int_69_103 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c104
+ bl_int_70_104 bl_int_69_104 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c105
+ bl_int_70_105 bl_int_69_105 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c106
+ bl_int_70_106 bl_int_69_106 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c107
+ bl_int_70_107 bl_int_69_107 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c108
+ bl_int_70_108 bl_int_69_108 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c109
+ bl_int_70_109 bl_int_69_109 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c110
+ bl_int_70_110 bl_int_69_110 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c111
+ bl_int_70_111 bl_int_69_111 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c112
+ bl_int_70_112 bl_int_69_112 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c113
+ bl_int_70_113 bl_int_69_113 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c114
+ bl_int_70_114 bl_int_69_114 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c115
+ bl_int_70_115 bl_int_69_115 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c116
+ bl_int_70_116 bl_int_69_116 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c117
+ bl_int_70_117 bl_int_69_117 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c118
+ bl_int_70_118 bl_int_69_118 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c119
+ bl_int_70_119 bl_int_69_119 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c120
+ bl_int_70_120 bl_int_69_120 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c121
+ bl_int_70_121 bl_int_69_121 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c122
+ bl_int_70_122 bl_int_69_122 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c123
+ bl_int_70_123 bl_int_69_123 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c124
+ bl_int_70_124 bl_int_69_124 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c125
+ bl_int_70_125 bl_int_69_125 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c126
+ bl_int_70_126 bl_int_69_126 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c127
+ bl_int_70_127 bl_int_69_127 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c128
+ bl_int_70_128 bl_int_69_128 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c129
+ bl_int_70_129 bl_int_69_129 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c130
+ bl_int_70_130 bl_int_69_130 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c131
+ bl_int_70_131 bl_int_69_131 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c132
+ bl_int_70_132 bl_int_69_132 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c133
+ bl_int_70_133 bl_int_69_133 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c134
+ bl_int_70_134 bl_int_69_134 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c135
+ bl_int_70_135 bl_int_69_135 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c136
+ bl_int_70_136 bl_int_69_136 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c137
+ bl_int_70_137 bl_int_69_137 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c138
+ bl_int_70_138 bl_int_69_138 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c139
+ bl_int_70_139 bl_int_69_139 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c140
+ bl_int_70_140 bl_int_69_140 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c141
+ bl_int_70_141 bl_int_69_141 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c142
+ bl_int_70_142 bl_int_69_142 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c143
+ bl_int_70_143 bl_int_69_143 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c144
+ bl_int_70_144 bl_int_69_144 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c145
+ bl_int_70_145 bl_int_69_145 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c146
+ bl_int_70_146 bl_int_69_146 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c147
+ bl_int_70_147 bl_int_69_147 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c148
+ bl_int_70_148 bl_int_69_148 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c149
+ bl_int_70_149 bl_int_69_149 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c150
+ bl_int_70_150 bl_int_69_150 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c151
+ bl_int_70_151 bl_int_69_151 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c152
+ bl_int_70_152 bl_int_69_152 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c153
+ bl_int_70_153 bl_int_69_153 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c154
+ bl_int_70_154 bl_int_69_154 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c155
+ bl_int_70_155 bl_int_69_155 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c156
+ bl_int_70_156 bl_int_69_156 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c157
+ bl_int_70_157 bl_int_69_157 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c158
+ bl_int_70_158 bl_int_69_158 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c159
+ bl_int_70_159 bl_int_69_159 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c160
+ bl_int_70_160 bl_int_69_160 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c161
+ bl_int_70_161 bl_int_69_161 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c162
+ bl_int_70_162 bl_int_69_162 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c163
+ bl_int_70_163 bl_int_69_163 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c164
+ bl_int_70_164 bl_int_69_164 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c165
+ bl_int_70_165 bl_int_69_165 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c166
+ bl_int_70_166 bl_int_69_166 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c167
+ bl_int_70_167 bl_int_69_167 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c168
+ bl_int_70_168 bl_int_69_168 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c169
+ bl_int_70_169 bl_int_69_169 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c170
+ bl_int_70_170 bl_int_69_170 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c171
+ bl_int_70_171 bl_int_69_171 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c172
+ bl_int_70_172 bl_int_69_172 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c173
+ bl_int_70_173 bl_int_69_173 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c174
+ bl_int_70_174 bl_int_69_174 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c175
+ bl_int_70_175 bl_int_69_175 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c176
+ bl_int_70_176 bl_int_69_176 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c177
+ bl_int_70_177 bl_int_69_177 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c178
+ bl_int_70_178 bl_int_69_178 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c179
+ bl_int_70_179 bl_int_69_179 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c180
+ bl_int_70_180 bl_int_69_180 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c181
+ bl_int_70_181 bl_int_69_181 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c182
+ bl_int_70_182 bl_int_69_182 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r70_c183
+ bl_int_70_183 bl_int_69_183 wl_0_70 gnd
+ sram_rom_base_one_cell
Xbit_r71_c0
+ bl_int_71_0 bl_int_70_0 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c1
+ bl_int_71_1 bl_int_70_1 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c2
+ bl_int_71_2 bl_int_70_2 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c3
+ bl_int_71_3 bl_int_70_3 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c4
+ bl_int_71_4 bl_int_70_4 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c5
+ bl_int_71_5 bl_int_70_5 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c6
+ bl_int_71_6 bl_int_70_6 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c7
+ bl_int_71_7 bl_int_70_7 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c8
+ bl_int_71_8 bl_int_70_8 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c9
+ bl_int_71_9 bl_int_70_9 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c10
+ bl_int_71_10 bl_int_70_10 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c11
+ bl_int_71_11 bl_int_70_11 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c12
+ bl_int_71_12 bl_int_70_12 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c13
+ bl_int_71_13 bl_int_70_13 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c14
+ bl_int_71_14 bl_int_70_14 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c15
+ bl_int_71_15 bl_int_70_15 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c16
+ bl_int_71_16 bl_int_70_16 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c17
+ bl_int_71_17 bl_int_70_17 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c18
+ bl_int_71_18 bl_int_70_18 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c19
+ bl_int_71_19 bl_int_70_19 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c20
+ bl_int_71_20 bl_int_70_20 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c21
+ bl_int_71_21 bl_int_70_21 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c22
+ bl_int_71_22 bl_int_70_22 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c23
+ bl_int_71_23 bl_int_70_23 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c24
+ bl_int_71_24 bl_int_70_24 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c25
+ bl_int_71_25 bl_int_70_25 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c26
+ bl_int_71_26 bl_int_70_26 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c27
+ bl_int_71_27 bl_int_70_27 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c28
+ bl_int_71_28 bl_int_70_28 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c29
+ bl_int_71_29 bl_int_70_29 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c30
+ bl_int_71_30 bl_int_70_30 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c31
+ bl_int_71_31 bl_int_70_31 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c32
+ bl_int_71_32 bl_int_70_32 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c33
+ bl_int_71_33 bl_int_70_33 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c34
+ bl_int_71_34 bl_int_70_34 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c35
+ bl_int_71_35 bl_int_70_35 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c36
+ bl_int_71_36 bl_int_70_36 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c37
+ bl_int_71_37 bl_int_70_37 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c38
+ bl_int_71_38 bl_int_70_38 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c39
+ bl_int_71_39 bl_int_70_39 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c40
+ bl_int_71_40 bl_int_70_40 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c41
+ bl_int_71_41 bl_int_70_41 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c42
+ bl_int_71_42 bl_int_70_42 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c43
+ bl_int_71_43 bl_int_70_43 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c44
+ bl_int_71_44 bl_int_70_44 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c45
+ bl_int_71_45 bl_int_70_45 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c46
+ bl_int_71_46 bl_int_70_46 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c47
+ bl_int_71_47 bl_int_70_47 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c48
+ bl_int_71_48 bl_int_70_48 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c49
+ bl_int_71_49 bl_int_70_49 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c50
+ bl_int_71_50 bl_int_70_50 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c51
+ bl_int_71_51 bl_int_70_51 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c52
+ bl_int_71_52 bl_int_70_52 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c53
+ bl_int_71_53 bl_int_70_53 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c54
+ bl_int_71_54 bl_int_70_54 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c55
+ bl_int_71_55 bl_int_70_55 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c56
+ bl_int_71_56 bl_int_70_56 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c57
+ bl_int_71_57 bl_int_70_57 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c58
+ bl_int_71_58 bl_int_70_58 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c59
+ bl_int_71_59 bl_int_70_59 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c60
+ bl_int_71_60 bl_int_70_60 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c61
+ bl_int_71_61 bl_int_70_61 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c62
+ bl_int_71_62 bl_int_70_62 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c63
+ bl_int_71_63 bl_int_70_63 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c64
+ bl_int_71_64 bl_int_70_64 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c65
+ bl_int_71_65 bl_int_70_65 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c66
+ bl_int_71_66 bl_int_70_66 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c67
+ bl_int_71_67 bl_int_70_67 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c68
+ bl_int_71_68 bl_int_70_68 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c69
+ bl_int_71_69 bl_int_70_69 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c70
+ bl_int_71_70 bl_int_70_70 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c71
+ bl_int_71_71 bl_int_70_71 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c72
+ bl_int_71_72 bl_int_70_72 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c73
+ bl_int_71_73 bl_int_70_73 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c74
+ bl_int_71_74 bl_int_70_74 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c75
+ bl_int_71_75 bl_int_70_75 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c76
+ bl_int_71_76 bl_int_70_76 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c77
+ bl_int_71_77 bl_int_70_77 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c78
+ bl_int_71_78 bl_int_70_78 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c79
+ bl_int_71_79 bl_int_70_79 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c80
+ bl_int_71_80 bl_int_70_80 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c81
+ bl_int_71_81 bl_int_70_81 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c82
+ bl_int_71_82 bl_int_70_82 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c83
+ bl_int_71_83 bl_int_70_83 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c84
+ bl_int_71_84 bl_int_70_84 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c85
+ bl_int_71_85 bl_int_70_85 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c86
+ bl_int_71_86 bl_int_70_86 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c87
+ bl_int_71_87 bl_int_70_87 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c88
+ bl_int_71_88 bl_int_70_88 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c89
+ bl_int_71_89 bl_int_70_89 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c90
+ bl_int_71_90 bl_int_70_90 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c91
+ bl_int_71_91 bl_int_70_91 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c92
+ bl_int_71_92 bl_int_70_92 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c93
+ bl_int_71_93 bl_int_70_93 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c94
+ bl_int_71_94 bl_int_70_94 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c95
+ bl_int_71_95 bl_int_70_95 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c96
+ bl_int_71_96 bl_int_70_96 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c97
+ bl_int_71_97 bl_int_70_97 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c98
+ bl_int_71_98 bl_int_70_98 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c99
+ bl_int_71_99 bl_int_70_99 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c100
+ bl_int_71_100 bl_int_70_100 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c101
+ bl_int_71_101 bl_int_70_101 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c102
+ bl_int_71_102 bl_int_70_102 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c103
+ bl_int_71_103 bl_int_70_103 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c104
+ bl_int_71_104 bl_int_70_104 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c105
+ bl_int_71_105 bl_int_70_105 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c106
+ bl_int_71_106 bl_int_70_106 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c107
+ bl_int_71_107 bl_int_70_107 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c108
+ bl_int_71_108 bl_int_70_108 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c109
+ bl_int_71_109 bl_int_70_109 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c110
+ bl_int_71_110 bl_int_70_110 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c111
+ bl_int_71_111 bl_int_70_111 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c112
+ bl_int_71_112 bl_int_70_112 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c113
+ bl_int_71_113 bl_int_70_113 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c114
+ bl_int_71_114 bl_int_70_114 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c115
+ bl_int_71_115 bl_int_70_115 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c116
+ bl_int_71_116 bl_int_70_116 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c117
+ bl_int_71_117 bl_int_70_117 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c118
+ bl_int_71_118 bl_int_70_118 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c119
+ bl_int_71_119 bl_int_70_119 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c120
+ bl_int_71_120 bl_int_70_120 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c121
+ bl_int_71_121 bl_int_70_121 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c122
+ bl_int_71_122 bl_int_70_122 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c123
+ bl_int_71_123 bl_int_70_123 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c124
+ bl_int_71_124 bl_int_70_124 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c125
+ bl_int_71_125 bl_int_70_125 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c126
+ bl_int_71_126 bl_int_70_126 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c127
+ bl_int_71_127 bl_int_70_127 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c128
+ bl_int_71_128 bl_int_70_128 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c129
+ bl_int_71_129 bl_int_70_129 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c130
+ bl_int_71_130 bl_int_70_130 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c131
+ bl_int_71_131 bl_int_70_131 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c132
+ bl_int_71_132 bl_int_70_132 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c133
+ bl_int_71_133 bl_int_70_133 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c134
+ bl_int_71_134 bl_int_70_134 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c135
+ bl_int_71_135 bl_int_70_135 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c136
+ bl_int_71_136 bl_int_70_136 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c137
+ bl_int_71_137 bl_int_70_137 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c138
+ bl_int_71_138 bl_int_70_138 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c139
+ bl_int_71_139 bl_int_70_139 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c140
+ bl_int_71_140 bl_int_70_140 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c141
+ bl_int_71_141 bl_int_70_141 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c142
+ bl_int_71_142 bl_int_70_142 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c143
+ bl_int_71_143 bl_int_70_143 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c144
+ bl_int_71_144 bl_int_70_144 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c145
+ bl_int_71_145 bl_int_70_145 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c146
+ bl_int_71_146 bl_int_70_146 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c147
+ bl_int_71_147 bl_int_70_147 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c148
+ bl_int_71_148 bl_int_70_148 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c149
+ bl_int_71_149 bl_int_70_149 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c150
+ bl_int_71_150 bl_int_70_150 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c151
+ bl_int_71_151 bl_int_70_151 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c152
+ bl_int_71_152 bl_int_70_152 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c153
+ bl_int_71_153 bl_int_70_153 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c154
+ bl_int_71_154 bl_int_70_154 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c155
+ bl_int_71_155 bl_int_70_155 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c156
+ bl_int_71_156 bl_int_70_156 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c157
+ bl_int_71_157 bl_int_70_157 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c158
+ bl_int_71_158 bl_int_70_158 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c159
+ bl_int_71_159 bl_int_70_159 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c160
+ bl_int_71_160 bl_int_70_160 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c161
+ bl_int_71_161 bl_int_70_161 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c162
+ bl_int_71_162 bl_int_70_162 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c163
+ bl_int_71_163 bl_int_70_163 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c164
+ bl_int_71_164 bl_int_70_164 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c165
+ bl_int_71_165 bl_int_70_165 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c166
+ bl_int_71_166 bl_int_70_166 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c167
+ bl_int_71_167 bl_int_70_167 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c168
+ bl_int_71_168 bl_int_70_168 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c169
+ bl_int_71_169 bl_int_70_169 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c170
+ bl_int_71_170 bl_int_70_170 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c171
+ bl_int_71_171 bl_int_70_171 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c172
+ bl_int_71_172 bl_int_70_172 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c173
+ bl_int_71_173 bl_int_70_173 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c174
+ bl_int_71_174 bl_int_70_174 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c175
+ bl_int_71_175 bl_int_70_175 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c176
+ bl_int_71_176 bl_int_70_176 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c177
+ bl_int_71_177 bl_int_70_177 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c178
+ bl_int_71_178 bl_int_70_178 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c179
+ bl_int_71_179 bl_int_70_179 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c180
+ bl_int_71_180 bl_int_70_180 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c181
+ bl_int_71_181 bl_int_70_181 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c182
+ bl_int_71_182 bl_int_70_182 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r71_c183
+ bl_int_71_183 bl_int_70_183 wl_0_71 gnd
+ sram_rom_base_one_cell
Xbit_r72_c0
+ bl_int_72_0 bl_int_71_0 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c1
+ bl_int_72_1 bl_int_71_1 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c2
+ bl_int_72_2 bl_int_71_2 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c3
+ bl_int_72_3 bl_int_71_3 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c4
+ bl_int_72_4 bl_int_71_4 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c5
+ bl_int_72_5 bl_int_71_5 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c6
+ bl_int_72_6 bl_int_71_6 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c7
+ bl_int_72_7 bl_int_71_7 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c8
+ bl_int_72_8 bl_int_71_8 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c9
+ bl_int_72_9 bl_int_71_9 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c10
+ bl_int_72_10 bl_int_71_10 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c11
+ bl_int_72_11 bl_int_71_11 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c12
+ bl_int_72_12 bl_int_71_12 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c13
+ bl_int_72_13 bl_int_71_13 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c14
+ bl_int_72_14 bl_int_71_14 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c15
+ bl_int_72_15 bl_int_71_15 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c16
+ bl_int_72_16 bl_int_71_16 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c17
+ bl_int_72_17 bl_int_71_17 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c18
+ bl_int_72_18 bl_int_71_18 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c19
+ bl_int_72_19 bl_int_71_19 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c20
+ bl_int_72_20 bl_int_71_20 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c21
+ bl_int_72_21 bl_int_71_21 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c22
+ bl_int_72_22 bl_int_71_22 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c23
+ bl_int_72_23 bl_int_71_23 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c24
+ bl_int_72_24 bl_int_71_24 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c25
+ bl_int_72_25 bl_int_71_25 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c26
+ bl_int_72_26 bl_int_71_26 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c27
+ bl_int_72_27 bl_int_71_27 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c28
+ bl_int_72_28 bl_int_71_28 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c29
+ bl_int_72_29 bl_int_71_29 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c30
+ bl_int_72_30 bl_int_71_30 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c31
+ bl_int_72_31 bl_int_71_31 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c32
+ bl_int_72_32 bl_int_71_32 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c33
+ bl_int_72_33 bl_int_71_33 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c34
+ bl_int_72_34 bl_int_71_34 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c35
+ bl_int_72_35 bl_int_71_35 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c36
+ bl_int_72_36 bl_int_71_36 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c37
+ bl_int_72_37 bl_int_71_37 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c38
+ bl_int_72_38 bl_int_71_38 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c39
+ bl_int_72_39 bl_int_71_39 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c40
+ bl_int_72_40 bl_int_71_40 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c41
+ bl_int_72_41 bl_int_71_41 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c42
+ bl_int_72_42 bl_int_71_42 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c43
+ bl_int_72_43 bl_int_71_43 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c44
+ bl_int_72_44 bl_int_71_44 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c45
+ bl_int_72_45 bl_int_71_45 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c46
+ bl_int_72_46 bl_int_71_46 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c47
+ bl_int_72_47 bl_int_71_47 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c48
+ bl_int_72_48 bl_int_71_48 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c49
+ bl_int_72_49 bl_int_71_49 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c50
+ bl_int_72_50 bl_int_71_50 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c51
+ bl_int_72_51 bl_int_71_51 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c52
+ bl_int_72_52 bl_int_71_52 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c53
+ bl_int_72_53 bl_int_71_53 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c54
+ bl_int_72_54 bl_int_71_54 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c55
+ bl_int_72_55 bl_int_71_55 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c56
+ bl_int_72_56 bl_int_71_56 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c57
+ bl_int_72_57 bl_int_71_57 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c58
+ bl_int_72_58 bl_int_71_58 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c59
+ bl_int_72_59 bl_int_71_59 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c60
+ bl_int_72_60 bl_int_71_60 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c61
+ bl_int_72_61 bl_int_71_61 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c62
+ bl_int_72_62 bl_int_71_62 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c63
+ bl_int_72_63 bl_int_71_63 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c64
+ bl_int_72_64 bl_int_71_64 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c65
+ bl_int_72_65 bl_int_71_65 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c66
+ bl_int_72_66 bl_int_71_66 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c67
+ bl_int_72_67 bl_int_71_67 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c68
+ bl_int_72_68 bl_int_71_68 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c69
+ bl_int_72_69 bl_int_71_69 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c70
+ bl_int_72_70 bl_int_71_70 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c71
+ bl_int_72_71 bl_int_71_71 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c72
+ bl_int_72_72 bl_int_71_72 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c73
+ bl_int_72_73 bl_int_71_73 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c74
+ bl_int_72_74 bl_int_71_74 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c75
+ bl_int_72_75 bl_int_71_75 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c76
+ bl_int_72_76 bl_int_71_76 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c77
+ bl_int_72_77 bl_int_71_77 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c78
+ bl_int_72_78 bl_int_71_78 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c79
+ bl_int_72_79 bl_int_71_79 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c80
+ bl_int_72_80 bl_int_71_80 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c81
+ bl_int_72_81 bl_int_71_81 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c82
+ bl_int_72_82 bl_int_71_82 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c83
+ bl_int_72_83 bl_int_71_83 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c84
+ bl_int_72_84 bl_int_71_84 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c85
+ bl_int_72_85 bl_int_71_85 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c86
+ bl_int_72_86 bl_int_71_86 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c87
+ bl_int_72_87 bl_int_71_87 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c88
+ bl_int_72_88 bl_int_71_88 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c89
+ bl_int_72_89 bl_int_71_89 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c90
+ bl_int_72_90 bl_int_71_90 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c91
+ bl_int_72_91 bl_int_71_91 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c92
+ bl_int_72_92 bl_int_71_92 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c93
+ bl_int_72_93 bl_int_71_93 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c94
+ bl_int_72_94 bl_int_71_94 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c95
+ bl_int_72_95 bl_int_71_95 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c96
+ bl_int_72_96 bl_int_71_96 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c97
+ bl_int_72_97 bl_int_71_97 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c98
+ bl_int_72_98 bl_int_71_98 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c99
+ bl_int_72_99 bl_int_71_99 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c100
+ bl_int_72_100 bl_int_71_100 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c101
+ bl_int_72_101 bl_int_71_101 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c102
+ bl_int_72_102 bl_int_71_102 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c103
+ bl_int_72_103 bl_int_71_103 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c104
+ bl_int_72_104 bl_int_71_104 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c105
+ bl_int_72_105 bl_int_71_105 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c106
+ bl_int_72_106 bl_int_71_106 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c107
+ bl_int_72_107 bl_int_71_107 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c108
+ bl_int_72_108 bl_int_71_108 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c109
+ bl_int_72_109 bl_int_71_109 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c110
+ bl_int_72_110 bl_int_71_110 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c111
+ bl_int_72_111 bl_int_71_111 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c112
+ bl_int_72_112 bl_int_71_112 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c113
+ bl_int_72_113 bl_int_71_113 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c114
+ bl_int_72_114 bl_int_71_114 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c115
+ bl_int_72_115 bl_int_71_115 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c116
+ bl_int_72_116 bl_int_71_116 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c117
+ bl_int_72_117 bl_int_71_117 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c118
+ bl_int_72_118 bl_int_71_118 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c119
+ bl_int_72_119 bl_int_71_119 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c120
+ bl_int_72_120 bl_int_71_120 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c121
+ bl_int_72_121 bl_int_71_121 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c122
+ bl_int_72_122 bl_int_71_122 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c123
+ bl_int_72_123 bl_int_71_123 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c124
+ bl_int_72_124 bl_int_71_124 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c125
+ bl_int_72_125 bl_int_71_125 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c126
+ bl_int_72_126 bl_int_71_126 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c127
+ bl_int_72_127 bl_int_71_127 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c128
+ bl_int_72_128 bl_int_71_128 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c129
+ bl_int_72_129 bl_int_71_129 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c130
+ bl_int_72_130 bl_int_71_130 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c131
+ bl_int_72_131 bl_int_71_131 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c132
+ bl_int_72_132 bl_int_71_132 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c133
+ bl_int_72_133 bl_int_71_133 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c134
+ bl_int_72_134 bl_int_71_134 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c135
+ bl_int_72_135 bl_int_71_135 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c136
+ bl_int_72_136 bl_int_71_136 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c137
+ bl_int_72_137 bl_int_71_137 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c138
+ bl_int_72_138 bl_int_71_138 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c139
+ bl_int_72_139 bl_int_71_139 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c140
+ bl_int_72_140 bl_int_71_140 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c141
+ bl_int_72_141 bl_int_71_141 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c142
+ bl_int_72_142 bl_int_71_142 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c143
+ bl_int_72_143 bl_int_71_143 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c144
+ bl_int_72_144 bl_int_71_144 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c145
+ bl_int_72_145 bl_int_71_145 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c146
+ bl_int_72_146 bl_int_71_146 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c147
+ bl_int_72_147 bl_int_71_147 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c148
+ bl_int_72_148 bl_int_71_148 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c149
+ bl_int_72_149 bl_int_71_149 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c150
+ bl_int_72_150 bl_int_71_150 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c151
+ bl_int_72_151 bl_int_71_151 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c152
+ bl_int_72_152 bl_int_71_152 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c153
+ bl_int_72_153 bl_int_71_153 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c154
+ bl_int_72_154 bl_int_71_154 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c155
+ bl_int_72_155 bl_int_71_155 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c156
+ bl_int_72_156 bl_int_71_156 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c157
+ bl_int_72_157 bl_int_71_157 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c158
+ bl_int_72_158 bl_int_71_158 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c159
+ bl_int_72_159 bl_int_71_159 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c160
+ bl_int_72_160 bl_int_71_160 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c161
+ bl_int_72_161 bl_int_71_161 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c162
+ bl_int_72_162 bl_int_71_162 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c163
+ bl_int_72_163 bl_int_71_163 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c164
+ bl_int_72_164 bl_int_71_164 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c165
+ bl_int_72_165 bl_int_71_165 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c166
+ bl_int_72_166 bl_int_71_166 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c167
+ bl_int_72_167 bl_int_71_167 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c168
+ bl_int_72_168 bl_int_71_168 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c169
+ bl_int_72_169 bl_int_71_169 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c170
+ bl_int_72_170 bl_int_71_170 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c171
+ bl_int_72_171 bl_int_71_171 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c172
+ bl_int_72_172 bl_int_71_172 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c173
+ bl_int_72_173 bl_int_71_173 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c174
+ bl_int_72_174 bl_int_71_174 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c175
+ bl_int_72_175 bl_int_71_175 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c176
+ bl_int_72_176 bl_int_71_176 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c177
+ bl_int_72_177 bl_int_71_177 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c178
+ bl_int_72_178 bl_int_71_178 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c179
+ bl_int_72_179 bl_int_71_179 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c180
+ bl_int_72_180 bl_int_71_180 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c181
+ bl_int_72_181 bl_int_71_181 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c182
+ bl_int_72_182 bl_int_71_182 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r72_c183
+ bl_int_72_183 bl_int_71_183 wl_0_72 gnd
+ sram_rom_base_one_cell
Xbit_r73_c0
+ bl_int_73_0 bl_int_72_0 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c1
+ bl_int_73_1 bl_int_72_1 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c2
+ bl_int_73_2 bl_int_72_2 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c3
+ bl_int_73_3 bl_int_72_3 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c4
+ bl_int_73_4 bl_int_72_4 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c5
+ bl_int_73_5 bl_int_72_5 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c6
+ bl_int_73_6 bl_int_72_6 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c7
+ bl_int_73_7 bl_int_72_7 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c8
+ bl_int_73_8 bl_int_72_8 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c9
+ bl_int_73_9 bl_int_72_9 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c10
+ bl_int_73_10 bl_int_72_10 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c11
+ bl_int_73_11 bl_int_72_11 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c12
+ bl_int_73_12 bl_int_72_12 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c13
+ bl_int_73_13 bl_int_72_13 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c14
+ bl_int_73_14 bl_int_72_14 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c15
+ bl_int_73_15 bl_int_72_15 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c16
+ bl_int_73_16 bl_int_72_16 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c17
+ bl_int_73_17 bl_int_72_17 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c18
+ bl_int_73_18 bl_int_72_18 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c19
+ bl_int_73_19 bl_int_72_19 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c20
+ bl_int_73_20 bl_int_72_20 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c21
+ bl_int_73_21 bl_int_72_21 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c22
+ bl_int_73_22 bl_int_72_22 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c23
+ bl_int_73_23 bl_int_72_23 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c24
+ bl_int_73_24 bl_int_72_24 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c25
+ bl_int_73_25 bl_int_72_25 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c26
+ bl_int_73_26 bl_int_72_26 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c27
+ bl_int_73_27 bl_int_72_27 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c28
+ bl_int_73_28 bl_int_72_28 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c29
+ bl_int_73_29 bl_int_72_29 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c30
+ bl_int_73_30 bl_int_72_30 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c31
+ bl_int_73_31 bl_int_72_31 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c32
+ bl_int_73_32 bl_int_72_32 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c33
+ bl_int_73_33 bl_int_72_33 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c34
+ bl_int_73_34 bl_int_72_34 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c35
+ bl_int_73_35 bl_int_72_35 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c36
+ bl_int_73_36 bl_int_72_36 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c37
+ bl_int_73_37 bl_int_72_37 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c38
+ bl_int_73_38 bl_int_72_38 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c39
+ bl_int_73_39 bl_int_72_39 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c40
+ bl_int_73_40 bl_int_72_40 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c41
+ bl_int_73_41 bl_int_72_41 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c42
+ bl_int_73_42 bl_int_72_42 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c43
+ bl_int_73_43 bl_int_72_43 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c44
+ bl_int_73_44 bl_int_72_44 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c45
+ bl_int_73_45 bl_int_72_45 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c46
+ bl_int_73_46 bl_int_72_46 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c47
+ bl_int_73_47 bl_int_72_47 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c48
+ bl_int_73_48 bl_int_72_48 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c49
+ bl_int_73_49 bl_int_72_49 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c50
+ bl_int_73_50 bl_int_72_50 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c51
+ bl_int_73_51 bl_int_72_51 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c52
+ bl_int_73_52 bl_int_72_52 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c53
+ bl_int_73_53 bl_int_72_53 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c54
+ bl_int_73_54 bl_int_72_54 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c55
+ bl_int_73_55 bl_int_72_55 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c56
+ bl_int_73_56 bl_int_72_56 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c57
+ bl_int_73_57 bl_int_72_57 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c58
+ bl_int_73_58 bl_int_72_58 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c59
+ bl_int_73_59 bl_int_72_59 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c60
+ bl_int_73_60 bl_int_72_60 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c61
+ bl_int_73_61 bl_int_72_61 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c62
+ bl_int_73_62 bl_int_72_62 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c63
+ bl_int_73_63 bl_int_72_63 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c64
+ bl_int_73_64 bl_int_72_64 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c65
+ bl_int_73_65 bl_int_72_65 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c66
+ bl_int_73_66 bl_int_72_66 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c67
+ bl_int_73_67 bl_int_72_67 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c68
+ bl_int_73_68 bl_int_72_68 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c69
+ bl_int_73_69 bl_int_72_69 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c70
+ bl_int_73_70 bl_int_72_70 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c71
+ bl_int_73_71 bl_int_72_71 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c72
+ bl_int_73_72 bl_int_72_72 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c73
+ bl_int_73_73 bl_int_72_73 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c74
+ bl_int_73_74 bl_int_72_74 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c75
+ bl_int_73_75 bl_int_72_75 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c76
+ bl_int_73_76 bl_int_72_76 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c77
+ bl_int_73_77 bl_int_72_77 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c78
+ bl_int_73_78 bl_int_72_78 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c79
+ bl_int_73_79 bl_int_72_79 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c80
+ bl_int_73_80 bl_int_72_80 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c81
+ bl_int_73_81 bl_int_72_81 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c82
+ bl_int_73_82 bl_int_72_82 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c83
+ bl_int_73_83 bl_int_72_83 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c84
+ bl_int_73_84 bl_int_72_84 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c85
+ bl_int_73_85 bl_int_72_85 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c86
+ bl_int_73_86 bl_int_72_86 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c87
+ bl_int_73_87 bl_int_72_87 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c88
+ bl_int_73_88 bl_int_72_88 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c89
+ bl_int_73_89 bl_int_72_89 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c90
+ bl_int_73_90 bl_int_72_90 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c91
+ bl_int_73_91 bl_int_72_91 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c92
+ bl_int_73_92 bl_int_72_92 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c93
+ bl_int_73_93 bl_int_72_93 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c94
+ bl_int_73_94 bl_int_72_94 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c95
+ bl_int_73_95 bl_int_72_95 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c96
+ bl_int_73_96 bl_int_72_96 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c97
+ bl_int_73_97 bl_int_72_97 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c98
+ bl_int_73_98 bl_int_72_98 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c99
+ bl_int_73_99 bl_int_72_99 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c100
+ bl_int_73_100 bl_int_72_100 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c101
+ bl_int_73_101 bl_int_72_101 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c102
+ bl_int_73_102 bl_int_72_102 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c103
+ bl_int_73_103 bl_int_72_103 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c104
+ bl_int_73_104 bl_int_72_104 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c105
+ bl_int_73_105 bl_int_72_105 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c106
+ bl_int_73_106 bl_int_72_106 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c107
+ bl_int_73_107 bl_int_72_107 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c108
+ bl_int_73_108 bl_int_72_108 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c109
+ bl_int_73_109 bl_int_72_109 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c110
+ bl_int_73_110 bl_int_72_110 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c111
+ bl_int_73_111 bl_int_72_111 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c112
+ bl_int_73_112 bl_int_72_112 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c113
+ bl_int_73_113 bl_int_72_113 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c114
+ bl_int_73_114 bl_int_72_114 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c115
+ bl_int_73_115 bl_int_72_115 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c116
+ bl_int_73_116 bl_int_72_116 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c117
+ bl_int_73_117 bl_int_72_117 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c118
+ bl_int_73_118 bl_int_72_118 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c119
+ bl_int_73_119 bl_int_72_119 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c120
+ bl_int_73_120 bl_int_72_120 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c121
+ bl_int_73_121 bl_int_72_121 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c122
+ bl_int_73_122 bl_int_72_122 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c123
+ bl_int_73_123 bl_int_72_123 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c124
+ bl_int_73_124 bl_int_72_124 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c125
+ bl_int_73_125 bl_int_72_125 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c126
+ bl_int_73_126 bl_int_72_126 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c127
+ bl_int_73_127 bl_int_72_127 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c128
+ bl_int_73_128 bl_int_72_128 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c129
+ bl_int_73_129 bl_int_72_129 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c130
+ bl_int_73_130 bl_int_72_130 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c131
+ bl_int_73_131 bl_int_72_131 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c132
+ bl_int_73_132 bl_int_72_132 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c133
+ bl_int_73_133 bl_int_72_133 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c134
+ bl_int_73_134 bl_int_72_134 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c135
+ bl_int_73_135 bl_int_72_135 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c136
+ bl_int_73_136 bl_int_72_136 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c137
+ bl_int_73_137 bl_int_72_137 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c138
+ bl_int_73_138 bl_int_72_138 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c139
+ bl_int_73_139 bl_int_72_139 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c140
+ bl_int_73_140 bl_int_72_140 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c141
+ bl_int_73_141 bl_int_72_141 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c142
+ bl_int_73_142 bl_int_72_142 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c143
+ bl_int_73_143 bl_int_72_143 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c144
+ bl_int_73_144 bl_int_72_144 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c145
+ bl_int_73_145 bl_int_72_145 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c146
+ bl_int_73_146 bl_int_72_146 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c147
+ bl_int_73_147 bl_int_72_147 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c148
+ bl_int_73_148 bl_int_72_148 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c149
+ bl_int_73_149 bl_int_72_149 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c150
+ bl_int_73_150 bl_int_72_150 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c151
+ bl_int_73_151 bl_int_72_151 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c152
+ bl_int_73_152 bl_int_72_152 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c153
+ bl_int_73_153 bl_int_72_153 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c154
+ bl_int_73_154 bl_int_72_154 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c155
+ bl_int_73_155 bl_int_72_155 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c156
+ bl_int_73_156 bl_int_72_156 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c157
+ bl_int_73_157 bl_int_72_157 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c158
+ bl_int_73_158 bl_int_72_158 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c159
+ bl_int_73_159 bl_int_72_159 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c160
+ bl_int_73_160 bl_int_72_160 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c161
+ bl_int_73_161 bl_int_72_161 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c162
+ bl_int_73_162 bl_int_72_162 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c163
+ bl_int_73_163 bl_int_72_163 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c164
+ bl_int_73_164 bl_int_72_164 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c165
+ bl_int_73_165 bl_int_72_165 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c166
+ bl_int_73_166 bl_int_72_166 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c167
+ bl_int_73_167 bl_int_72_167 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c168
+ bl_int_73_168 bl_int_72_168 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c169
+ bl_int_73_169 bl_int_72_169 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c170
+ bl_int_73_170 bl_int_72_170 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c171
+ bl_int_73_171 bl_int_72_171 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c172
+ bl_int_73_172 bl_int_72_172 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c173
+ bl_int_73_173 bl_int_72_173 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c174
+ bl_int_73_174 bl_int_72_174 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c175
+ bl_int_73_175 bl_int_72_175 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c176
+ bl_int_73_176 bl_int_72_176 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c177
+ bl_int_73_177 bl_int_72_177 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c178
+ bl_int_73_178 bl_int_72_178 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c179
+ bl_int_73_179 bl_int_72_179 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c180
+ bl_int_73_180 bl_int_72_180 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c181
+ bl_int_73_181 bl_int_72_181 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c182
+ bl_int_73_182 bl_int_72_182 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r73_c183
+ bl_int_73_183 bl_int_72_183 wl_0_73 gnd
+ sram_rom_base_one_cell
Xbit_r74_c0
+ bl_int_74_0 bl_int_73_0 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c1
+ bl_int_74_1 bl_int_73_1 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c2
+ bl_int_74_2 bl_int_73_2 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c3
+ bl_int_74_3 bl_int_73_3 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c4
+ bl_int_74_4 bl_int_73_4 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c5
+ bl_int_74_5 bl_int_73_5 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c6
+ bl_int_74_6 bl_int_73_6 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c7
+ bl_int_74_7 bl_int_73_7 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c8
+ bl_int_74_8 bl_int_73_8 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c9
+ bl_int_74_9 bl_int_73_9 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c10
+ bl_int_74_10 bl_int_73_10 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c11
+ bl_int_74_11 bl_int_73_11 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c12
+ bl_int_74_12 bl_int_73_12 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c13
+ bl_int_74_13 bl_int_73_13 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c14
+ bl_int_74_14 bl_int_73_14 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c15
+ bl_int_74_15 bl_int_73_15 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c16
+ bl_int_74_16 bl_int_73_16 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c17
+ bl_int_74_17 bl_int_73_17 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c18
+ bl_int_74_18 bl_int_73_18 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c19
+ bl_int_74_19 bl_int_73_19 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c20
+ bl_int_74_20 bl_int_73_20 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c21
+ bl_int_74_21 bl_int_73_21 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c22
+ bl_int_74_22 bl_int_73_22 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c23
+ bl_int_74_23 bl_int_73_23 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c24
+ bl_int_74_24 bl_int_73_24 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c25
+ bl_int_74_25 bl_int_73_25 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c26
+ bl_int_74_26 bl_int_73_26 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c27
+ bl_int_74_27 bl_int_73_27 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c28
+ bl_int_74_28 bl_int_73_28 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c29
+ bl_int_74_29 bl_int_73_29 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c30
+ bl_int_74_30 bl_int_73_30 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c31
+ bl_int_74_31 bl_int_73_31 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c32
+ bl_int_74_32 bl_int_73_32 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c33
+ bl_int_74_33 bl_int_73_33 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c34
+ bl_int_74_34 bl_int_73_34 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c35
+ bl_int_74_35 bl_int_73_35 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c36
+ bl_int_74_36 bl_int_73_36 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c37
+ bl_int_74_37 bl_int_73_37 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c38
+ bl_int_74_38 bl_int_73_38 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c39
+ bl_int_74_39 bl_int_73_39 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c40
+ bl_int_74_40 bl_int_73_40 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c41
+ bl_int_74_41 bl_int_73_41 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c42
+ bl_int_74_42 bl_int_73_42 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c43
+ bl_int_74_43 bl_int_73_43 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c44
+ bl_int_74_44 bl_int_73_44 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c45
+ bl_int_74_45 bl_int_73_45 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c46
+ bl_int_74_46 bl_int_73_46 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c47
+ bl_int_74_47 bl_int_73_47 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c48
+ bl_int_74_48 bl_int_73_48 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c49
+ bl_int_74_49 bl_int_73_49 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c50
+ bl_int_74_50 bl_int_73_50 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c51
+ bl_int_74_51 bl_int_73_51 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c52
+ bl_int_74_52 bl_int_73_52 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c53
+ bl_int_74_53 bl_int_73_53 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c54
+ bl_int_74_54 bl_int_73_54 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c55
+ bl_int_74_55 bl_int_73_55 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c56
+ bl_int_74_56 bl_int_73_56 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c57
+ bl_int_74_57 bl_int_73_57 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c58
+ bl_int_74_58 bl_int_73_58 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c59
+ bl_int_74_59 bl_int_73_59 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c60
+ bl_int_74_60 bl_int_73_60 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c61
+ bl_int_74_61 bl_int_73_61 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c62
+ bl_int_74_62 bl_int_73_62 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c63
+ bl_int_74_63 bl_int_73_63 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c64
+ bl_int_74_64 bl_int_73_64 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c65
+ bl_int_74_65 bl_int_73_65 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c66
+ bl_int_74_66 bl_int_73_66 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c67
+ bl_int_74_67 bl_int_73_67 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c68
+ bl_int_74_68 bl_int_73_68 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c69
+ bl_int_74_69 bl_int_73_69 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c70
+ bl_int_74_70 bl_int_73_70 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c71
+ bl_int_74_71 bl_int_73_71 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c72
+ bl_int_74_72 bl_int_73_72 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c73
+ bl_int_74_73 bl_int_73_73 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c74
+ bl_int_74_74 bl_int_73_74 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c75
+ bl_int_74_75 bl_int_73_75 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c76
+ bl_int_74_76 bl_int_73_76 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c77
+ bl_int_74_77 bl_int_73_77 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c78
+ bl_int_74_78 bl_int_73_78 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c79
+ bl_int_74_79 bl_int_73_79 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c80
+ bl_int_74_80 bl_int_73_80 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c81
+ bl_int_74_81 bl_int_73_81 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c82
+ bl_int_74_82 bl_int_73_82 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c83
+ bl_int_74_83 bl_int_73_83 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c84
+ bl_int_74_84 bl_int_73_84 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c85
+ bl_int_74_85 bl_int_73_85 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c86
+ bl_int_74_86 bl_int_73_86 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c87
+ bl_int_74_87 bl_int_73_87 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c88
+ bl_int_74_88 bl_int_73_88 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c89
+ bl_int_74_89 bl_int_73_89 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c90
+ bl_int_74_90 bl_int_73_90 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c91
+ bl_int_74_91 bl_int_73_91 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c92
+ bl_int_74_92 bl_int_73_92 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c93
+ bl_int_74_93 bl_int_73_93 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c94
+ bl_int_74_94 bl_int_73_94 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c95
+ bl_int_74_95 bl_int_73_95 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c96
+ bl_int_74_96 bl_int_73_96 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c97
+ bl_int_74_97 bl_int_73_97 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c98
+ bl_int_74_98 bl_int_73_98 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c99
+ bl_int_74_99 bl_int_73_99 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c100
+ bl_int_74_100 bl_int_73_100 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c101
+ bl_int_74_101 bl_int_73_101 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c102
+ bl_int_74_102 bl_int_73_102 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c103
+ bl_int_74_103 bl_int_73_103 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c104
+ bl_int_74_104 bl_int_73_104 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c105
+ bl_int_74_105 bl_int_73_105 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c106
+ bl_int_74_106 bl_int_73_106 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c107
+ bl_int_74_107 bl_int_73_107 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c108
+ bl_int_74_108 bl_int_73_108 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c109
+ bl_int_74_109 bl_int_73_109 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c110
+ bl_int_74_110 bl_int_73_110 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c111
+ bl_int_74_111 bl_int_73_111 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c112
+ bl_int_74_112 bl_int_73_112 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c113
+ bl_int_74_113 bl_int_73_113 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c114
+ bl_int_74_114 bl_int_73_114 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c115
+ bl_int_74_115 bl_int_73_115 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c116
+ bl_int_74_116 bl_int_73_116 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c117
+ bl_int_74_117 bl_int_73_117 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c118
+ bl_int_74_118 bl_int_73_118 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c119
+ bl_int_74_119 bl_int_73_119 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c120
+ bl_int_74_120 bl_int_73_120 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c121
+ bl_int_74_121 bl_int_73_121 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c122
+ bl_int_74_122 bl_int_73_122 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c123
+ bl_int_74_123 bl_int_73_123 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c124
+ bl_int_74_124 bl_int_73_124 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c125
+ bl_int_74_125 bl_int_73_125 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c126
+ bl_int_74_126 bl_int_73_126 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c127
+ bl_int_74_127 bl_int_73_127 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c128
+ bl_int_74_128 bl_int_73_128 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c129
+ bl_int_74_129 bl_int_73_129 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c130
+ bl_int_74_130 bl_int_73_130 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c131
+ bl_int_74_131 bl_int_73_131 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c132
+ bl_int_74_132 bl_int_73_132 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c133
+ bl_int_74_133 bl_int_73_133 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c134
+ bl_int_74_134 bl_int_73_134 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c135
+ bl_int_74_135 bl_int_73_135 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c136
+ bl_int_74_136 bl_int_73_136 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c137
+ bl_int_74_137 bl_int_73_137 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c138
+ bl_int_74_138 bl_int_73_138 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c139
+ bl_int_74_139 bl_int_73_139 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c140
+ bl_int_74_140 bl_int_73_140 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c141
+ bl_int_74_141 bl_int_73_141 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c142
+ bl_int_74_142 bl_int_73_142 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c143
+ bl_int_74_143 bl_int_73_143 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c144
+ bl_int_74_144 bl_int_73_144 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c145
+ bl_int_74_145 bl_int_73_145 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c146
+ bl_int_74_146 bl_int_73_146 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c147
+ bl_int_74_147 bl_int_73_147 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c148
+ bl_int_74_148 bl_int_73_148 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c149
+ bl_int_74_149 bl_int_73_149 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c150
+ bl_int_74_150 bl_int_73_150 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c151
+ bl_int_74_151 bl_int_73_151 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c152
+ bl_int_74_152 bl_int_73_152 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c153
+ bl_int_74_153 bl_int_73_153 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c154
+ bl_int_74_154 bl_int_73_154 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c155
+ bl_int_74_155 bl_int_73_155 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c156
+ bl_int_74_156 bl_int_73_156 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c157
+ bl_int_74_157 bl_int_73_157 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c158
+ bl_int_74_158 bl_int_73_158 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c159
+ bl_int_74_159 bl_int_73_159 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c160
+ bl_int_74_160 bl_int_73_160 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c161
+ bl_int_74_161 bl_int_73_161 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c162
+ bl_int_74_162 bl_int_73_162 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c163
+ bl_int_74_163 bl_int_73_163 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c164
+ bl_int_74_164 bl_int_73_164 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c165
+ bl_int_74_165 bl_int_73_165 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c166
+ bl_int_74_166 bl_int_73_166 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c167
+ bl_int_74_167 bl_int_73_167 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c168
+ bl_int_74_168 bl_int_73_168 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c169
+ bl_int_74_169 bl_int_73_169 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c170
+ bl_int_74_170 bl_int_73_170 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c171
+ bl_int_74_171 bl_int_73_171 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c172
+ bl_int_74_172 bl_int_73_172 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c173
+ bl_int_74_173 bl_int_73_173 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c174
+ bl_int_74_174 bl_int_73_174 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c175
+ bl_int_74_175 bl_int_73_175 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c176
+ bl_int_74_176 bl_int_73_176 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c177
+ bl_int_74_177 bl_int_73_177 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c178
+ bl_int_74_178 bl_int_73_178 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c179
+ bl_int_74_179 bl_int_73_179 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c180
+ bl_int_74_180 bl_int_73_180 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c181
+ bl_int_74_181 bl_int_73_181 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c182
+ bl_int_74_182 bl_int_73_182 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r74_c183
+ bl_int_74_183 bl_int_73_183 wl_0_74 gnd
+ sram_rom_base_one_cell
Xbit_r75_c0
+ bl_int_75_0 bl_int_74_0 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c1
+ bl_int_75_1 bl_int_74_1 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c2
+ bl_int_75_2 bl_int_74_2 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c3
+ bl_int_75_3 bl_int_74_3 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c4
+ bl_int_75_4 bl_int_74_4 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c5
+ bl_int_75_5 bl_int_74_5 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c6
+ bl_int_75_6 bl_int_74_6 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c7
+ bl_int_75_7 bl_int_74_7 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c8
+ bl_int_75_8 bl_int_74_8 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c9
+ bl_int_75_9 bl_int_74_9 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c10
+ bl_int_75_10 bl_int_74_10 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c11
+ bl_int_75_11 bl_int_74_11 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c12
+ bl_int_75_12 bl_int_74_12 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c13
+ bl_int_75_13 bl_int_74_13 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c14
+ bl_int_75_14 bl_int_74_14 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c15
+ bl_int_75_15 bl_int_74_15 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c16
+ bl_int_75_16 bl_int_74_16 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c17
+ bl_int_75_17 bl_int_74_17 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c18
+ bl_int_75_18 bl_int_74_18 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c19
+ bl_int_75_19 bl_int_74_19 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c20
+ bl_int_75_20 bl_int_74_20 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c21
+ bl_int_75_21 bl_int_74_21 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c22
+ bl_int_75_22 bl_int_74_22 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c23
+ bl_int_75_23 bl_int_74_23 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c24
+ bl_int_75_24 bl_int_74_24 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c25
+ bl_int_75_25 bl_int_74_25 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c26
+ bl_int_75_26 bl_int_74_26 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c27
+ bl_int_75_27 bl_int_74_27 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c28
+ bl_int_75_28 bl_int_74_28 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c29
+ bl_int_75_29 bl_int_74_29 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c30
+ bl_int_75_30 bl_int_74_30 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c31
+ bl_int_75_31 bl_int_74_31 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c32
+ bl_int_75_32 bl_int_74_32 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c33
+ bl_int_75_33 bl_int_74_33 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c34
+ bl_int_75_34 bl_int_74_34 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c35
+ bl_int_75_35 bl_int_74_35 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c36
+ bl_int_75_36 bl_int_74_36 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c37
+ bl_int_75_37 bl_int_74_37 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c38
+ bl_int_75_38 bl_int_74_38 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c39
+ bl_int_75_39 bl_int_74_39 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c40
+ bl_int_75_40 bl_int_74_40 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c41
+ bl_int_75_41 bl_int_74_41 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c42
+ bl_int_75_42 bl_int_74_42 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c43
+ bl_int_75_43 bl_int_74_43 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c44
+ bl_int_75_44 bl_int_74_44 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c45
+ bl_int_75_45 bl_int_74_45 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c46
+ bl_int_75_46 bl_int_74_46 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c47
+ bl_int_75_47 bl_int_74_47 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c48
+ bl_int_75_48 bl_int_74_48 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c49
+ bl_int_75_49 bl_int_74_49 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c50
+ bl_int_75_50 bl_int_74_50 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c51
+ bl_int_75_51 bl_int_74_51 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c52
+ bl_int_75_52 bl_int_74_52 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c53
+ bl_int_75_53 bl_int_74_53 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c54
+ bl_int_75_54 bl_int_74_54 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c55
+ bl_int_75_55 bl_int_74_55 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c56
+ bl_int_75_56 bl_int_74_56 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c57
+ bl_int_75_57 bl_int_74_57 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c58
+ bl_int_75_58 bl_int_74_58 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c59
+ bl_int_75_59 bl_int_74_59 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c60
+ bl_int_75_60 bl_int_74_60 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c61
+ bl_int_75_61 bl_int_74_61 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c62
+ bl_int_75_62 bl_int_74_62 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c63
+ bl_int_75_63 bl_int_74_63 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c64
+ bl_int_75_64 bl_int_74_64 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c65
+ bl_int_75_65 bl_int_74_65 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c66
+ bl_int_75_66 bl_int_74_66 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c67
+ bl_int_75_67 bl_int_74_67 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c68
+ bl_int_75_68 bl_int_74_68 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c69
+ bl_int_75_69 bl_int_74_69 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c70
+ bl_int_75_70 bl_int_74_70 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c71
+ bl_int_75_71 bl_int_74_71 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c72
+ bl_int_75_72 bl_int_74_72 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c73
+ bl_int_75_73 bl_int_74_73 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c74
+ bl_int_75_74 bl_int_74_74 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c75
+ bl_int_75_75 bl_int_74_75 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c76
+ bl_int_75_76 bl_int_74_76 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c77
+ bl_int_75_77 bl_int_74_77 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c78
+ bl_int_75_78 bl_int_74_78 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c79
+ bl_int_75_79 bl_int_74_79 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c80
+ bl_int_75_80 bl_int_74_80 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c81
+ bl_int_75_81 bl_int_74_81 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c82
+ bl_int_75_82 bl_int_74_82 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c83
+ bl_int_75_83 bl_int_74_83 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c84
+ bl_int_75_84 bl_int_74_84 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c85
+ bl_int_75_85 bl_int_74_85 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c86
+ bl_int_75_86 bl_int_74_86 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c87
+ bl_int_75_87 bl_int_74_87 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c88
+ bl_int_75_88 bl_int_74_88 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c89
+ bl_int_75_89 bl_int_74_89 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c90
+ bl_int_75_90 bl_int_74_90 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c91
+ bl_int_75_91 bl_int_74_91 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c92
+ bl_int_75_92 bl_int_74_92 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c93
+ bl_int_75_93 bl_int_74_93 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c94
+ bl_int_75_94 bl_int_74_94 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c95
+ bl_int_75_95 bl_int_74_95 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c96
+ bl_int_75_96 bl_int_74_96 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c97
+ bl_int_75_97 bl_int_74_97 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c98
+ bl_int_75_98 bl_int_74_98 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c99
+ bl_int_75_99 bl_int_74_99 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c100
+ bl_int_75_100 bl_int_74_100 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c101
+ bl_int_75_101 bl_int_74_101 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c102
+ bl_int_75_102 bl_int_74_102 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c103
+ bl_int_75_103 bl_int_74_103 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c104
+ bl_int_75_104 bl_int_74_104 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c105
+ bl_int_75_105 bl_int_74_105 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c106
+ bl_int_75_106 bl_int_74_106 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c107
+ bl_int_75_107 bl_int_74_107 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c108
+ bl_int_75_108 bl_int_74_108 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c109
+ bl_int_75_109 bl_int_74_109 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c110
+ bl_int_75_110 bl_int_74_110 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c111
+ bl_int_75_111 bl_int_74_111 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c112
+ bl_int_75_112 bl_int_74_112 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c113
+ bl_int_75_113 bl_int_74_113 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c114
+ bl_int_75_114 bl_int_74_114 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c115
+ bl_int_75_115 bl_int_74_115 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c116
+ bl_int_75_116 bl_int_74_116 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c117
+ bl_int_75_117 bl_int_74_117 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c118
+ bl_int_75_118 bl_int_74_118 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c119
+ bl_int_75_119 bl_int_74_119 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c120
+ bl_int_75_120 bl_int_74_120 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c121
+ bl_int_75_121 bl_int_74_121 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c122
+ bl_int_75_122 bl_int_74_122 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c123
+ bl_int_75_123 bl_int_74_123 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c124
+ bl_int_75_124 bl_int_74_124 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c125
+ bl_int_75_125 bl_int_74_125 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c126
+ bl_int_75_126 bl_int_74_126 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c127
+ bl_int_75_127 bl_int_74_127 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c128
+ bl_int_75_128 bl_int_74_128 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c129
+ bl_int_75_129 bl_int_74_129 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c130
+ bl_int_75_130 bl_int_74_130 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c131
+ bl_int_75_131 bl_int_74_131 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c132
+ bl_int_75_132 bl_int_74_132 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c133
+ bl_int_75_133 bl_int_74_133 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c134
+ bl_int_75_134 bl_int_74_134 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c135
+ bl_int_75_135 bl_int_74_135 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c136
+ bl_int_75_136 bl_int_74_136 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c137
+ bl_int_75_137 bl_int_74_137 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c138
+ bl_int_75_138 bl_int_74_138 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c139
+ bl_int_75_139 bl_int_74_139 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c140
+ bl_int_75_140 bl_int_74_140 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c141
+ bl_int_75_141 bl_int_74_141 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c142
+ bl_int_75_142 bl_int_74_142 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c143
+ bl_int_75_143 bl_int_74_143 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c144
+ bl_int_75_144 bl_int_74_144 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c145
+ bl_int_75_145 bl_int_74_145 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c146
+ bl_int_75_146 bl_int_74_146 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c147
+ bl_int_75_147 bl_int_74_147 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c148
+ bl_int_75_148 bl_int_74_148 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c149
+ bl_int_75_149 bl_int_74_149 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c150
+ bl_int_75_150 bl_int_74_150 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c151
+ bl_int_75_151 bl_int_74_151 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c152
+ bl_int_75_152 bl_int_74_152 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c153
+ bl_int_75_153 bl_int_74_153 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c154
+ bl_int_75_154 bl_int_74_154 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c155
+ bl_int_75_155 bl_int_74_155 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c156
+ bl_int_75_156 bl_int_74_156 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c157
+ bl_int_75_157 bl_int_74_157 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c158
+ bl_int_75_158 bl_int_74_158 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c159
+ bl_int_75_159 bl_int_74_159 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c160
+ bl_int_75_160 bl_int_74_160 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c161
+ bl_int_75_161 bl_int_74_161 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c162
+ bl_int_75_162 bl_int_74_162 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c163
+ bl_int_75_163 bl_int_74_163 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c164
+ bl_int_75_164 bl_int_74_164 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c165
+ bl_int_75_165 bl_int_74_165 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c166
+ bl_int_75_166 bl_int_74_166 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c167
+ bl_int_75_167 bl_int_74_167 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c168
+ bl_int_75_168 bl_int_74_168 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c169
+ bl_int_75_169 bl_int_74_169 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c170
+ bl_int_75_170 bl_int_74_170 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c171
+ bl_int_75_171 bl_int_74_171 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c172
+ bl_int_75_172 bl_int_74_172 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c173
+ bl_int_75_173 bl_int_74_173 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c174
+ bl_int_75_174 bl_int_74_174 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c175
+ bl_int_75_175 bl_int_74_175 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c176
+ bl_int_75_176 bl_int_74_176 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c177
+ bl_int_75_177 bl_int_74_177 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c178
+ bl_int_75_178 bl_int_74_178 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c179
+ bl_int_75_179 bl_int_74_179 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c180
+ bl_int_75_180 bl_int_74_180 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c181
+ bl_int_75_181 bl_int_74_181 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c182
+ bl_int_75_182 bl_int_74_182 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r75_c183
+ bl_int_75_183 bl_int_74_183 wl_0_75 gnd
+ sram_rom_base_one_cell
Xbit_r76_c0
+ bl_int_76_0 bl_int_75_0 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c1
+ bl_int_76_1 bl_int_75_1 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c2
+ bl_int_76_2 bl_int_75_2 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c3
+ bl_int_76_3 bl_int_75_3 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c4
+ bl_int_76_4 bl_int_75_4 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c5
+ bl_int_76_5 bl_int_75_5 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c6
+ bl_int_76_6 bl_int_75_6 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c7
+ bl_int_76_7 bl_int_75_7 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c8
+ bl_int_76_8 bl_int_75_8 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c9
+ bl_int_76_9 bl_int_75_9 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c10
+ bl_int_76_10 bl_int_75_10 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c11
+ bl_int_76_11 bl_int_75_11 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c12
+ bl_int_76_12 bl_int_75_12 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c13
+ bl_int_76_13 bl_int_75_13 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c14
+ bl_int_76_14 bl_int_75_14 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c15
+ bl_int_76_15 bl_int_75_15 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c16
+ bl_int_76_16 bl_int_75_16 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c17
+ bl_int_76_17 bl_int_75_17 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c18
+ bl_int_76_18 bl_int_75_18 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c19
+ bl_int_76_19 bl_int_75_19 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c20
+ bl_int_76_20 bl_int_75_20 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c21
+ bl_int_76_21 bl_int_75_21 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c22
+ bl_int_76_22 bl_int_75_22 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c23
+ bl_int_76_23 bl_int_75_23 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c24
+ bl_int_76_24 bl_int_75_24 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c25
+ bl_int_76_25 bl_int_75_25 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c26
+ bl_int_76_26 bl_int_75_26 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c27
+ bl_int_76_27 bl_int_75_27 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c28
+ bl_int_76_28 bl_int_75_28 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c29
+ bl_int_76_29 bl_int_75_29 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c30
+ bl_int_76_30 bl_int_75_30 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c31
+ bl_int_76_31 bl_int_75_31 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c32
+ bl_int_76_32 bl_int_75_32 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c33
+ bl_int_76_33 bl_int_75_33 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c34
+ bl_int_76_34 bl_int_75_34 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c35
+ bl_int_76_35 bl_int_75_35 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c36
+ bl_int_76_36 bl_int_75_36 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c37
+ bl_int_76_37 bl_int_75_37 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c38
+ bl_int_76_38 bl_int_75_38 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c39
+ bl_int_76_39 bl_int_75_39 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c40
+ bl_int_76_40 bl_int_75_40 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c41
+ bl_int_76_41 bl_int_75_41 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c42
+ bl_int_76_42 bl_int_75_42 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c43
+ bl_int_76_43 bl_int_75_43 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c44
+ bl_int_76_44 bl_int_75_44 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c45
+ bl_int_76_45 bl_int_75_45 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c46
+ bl_int_76_46 bl_int_75_46 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c47
+ bl_int_76_47 bl_int_75_47 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c48
+ bl_int_76_48 bl_int_75_48 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c49
+ bl_int_76_49 bl_int_75_49 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c50
+ bl_int_76_50 bl_int_75_50 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c51
+ bl_int_76_51 bl_int_75_51 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c52
+ bl_int_76_52 bl_int_75_52 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c53
+ bl_int_76_53 bl_int_75_53 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c54
+ bl_int_76_54 bl_int_75_54 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c55
+ bl_int_76_55 bl_int_75_55 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c56
+ bl_int_76_56 bl_int_75_56 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c57
+ bl_int_76_57 bl_int_75_57 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c58
+ bl_int_76_58 bl_int_75_58 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c59
+ bl_int_76_59 bl_int_75_59 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c60
+ bl_int_76_60 bl_int_75_60 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c61
+ bl_int_76_61 bl_int_75_61 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c62
+ bl_int_76_62 bl_int_75_62 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c63
+ bl_int_76_63 bl_int_75_63 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c64
+ bl_int_76_64 bl_int_75_64 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c65
+ bl_int_76_65 bl_int_75_65 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c66
+ bl_int_76_66 bl_int_75_66 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c67
+ bl_int_76_67 bl_int_75_67 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c68
+ bl_int_76_68 bl_int_75_68 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c69
+ bl_int_76_69 bl_int_75_69 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c70
+ bl_int_76_70 bl_int_75_70 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c71
+ bl_int_76_71 bl_int_75_71 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c72
+ bl_int_76_72 bl_int_75_72 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c73
+ bl_int_76_73 bl_int_75_73 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c74
+ bl_int_76_74 bl_int_75_74 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c75
+ bl_int_76_75 bl_int_75_75 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c76
+ bl_int_76_76 bl_int_75_76 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c77
+ bl_int_76_77 bl_int_75_77 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c78
+ bl_int_76_78 bl_int_75_78 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c79
+ bl_int_76_79 bl_int_75_79 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c80
+ bl_int_76_80 bl_int_75_80 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c81
+ bl_int_76_81 bl_int_75_81 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c82
+ bl_int_76_82 bl_int_75_82 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c83
+ bl_int_76_83 bl_int_75_83 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c84
+ bl_int_76_84 bl_int_75_84 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c85
+ bl_int_76_85 bl_int_75_85 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c86
+ bl_int_76_86 bl_int_75_86 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c87
+ bl_int_76_87 bl_int_75_87 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c88
+ bl_int_76_88 bl_int_75_88 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c89
+ bl_int_76_89 bl_int_75_89 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c90
+ bl_int_76_90 bl_int_75_90 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c91
+ bl_int_76_91 bl_int_75_91 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c92
+ bl_int_76_92 bl_int_75_92 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c93
+ bl_int_76_93 bl_int_75_93 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c94
+ bl_int_76_94 bl_int_75_94 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c95
+ bl_int_76_95 bl_int_75_95 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c96
+ bl_int_76_96 bl_int_75_96 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c97
+ bl_int_76_97 bl_int_75_97 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c98
+ bl_int_76_98 bl_int_75_98 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c99
+ bl_int_76_99 bl_int_75_99 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c100
+ bl_int_76_100 bl_int_75_100 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c101
+ bl_int_76_101 bl_int_75_101 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c102
+ bl_int_76_102 bl_int_75_102 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c103
+ bl_int_76_103 bl_int_75_103 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c104
+ bl_int_76_104 bl_int_75_104 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c105
+ bl_int_76_105 bl_int_75_105 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c106
+ bl_int_76_106 bl_int_75_106 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c107
+ bl_int_76_107 bl_int_75_107 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c108
+ bl_int_76_108 bl_int_75_108 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c109
+ bl_int_76_109 bl_int_75_109 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c110
+ bl_int_76_110 bl_int_75_110 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c111
+ bl_int_76_111 bl_int_75_111 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c112
+ bl_int_76_112 bl_int_75_112 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c113
+ bl_int_76_113 bl_int_75_113 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c114
+ bl_int_76_114 bl_int_75_114 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c115
+ bl_int_76_115 bl_int_75_115 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c116
+ bl_int_76_116 bl_int_75_116 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c117
+ bl_int_76_117 bl_int_75_117 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c118
+ bl_int_76_118 bl_int_75_118 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c119
+ bl_int_76_119 bl_int_75_119 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c120
+ bl_int_76_120 bl_int_75_120 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c121
+ bl_int_76_121 bl_int_75_121 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c122
+ bl_int_76_122 bl_int_75_122 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c123
+ bl_int_76_123 bl_int_75_123 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c124
+ bl_int_76_124 bl_int_75_124 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c125
+ bl_int_76_125 bl_int_75_125 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c126
+ bl_int_76_126 bl_int_75_126 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c127
+ bl_int_76_127 bl_int_75_127 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c128
+ bl_int_76_128 bl_int_75_128 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c129
+ bl_int_76_129 bl_int_75_129 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c130
+ bl_int_76_130 bl_int_75_130 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c131
+ bl_int_76_131 bl_int_75_131 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c132
+ bl_int_76_132 bl_int_75_132 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c133
+ bl_int_76_133 bl_int_75_133 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c134
+ bl_int_76_134 bl_int_75_134 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c135
+ bl_int_76_135 bl_int_75_135 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c136
+ bl_int_76_136 bl_int_75_136 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c137
+ bl_int_76_137 bl_int_75_137 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c138
+ bl_int_76_138 bl_int_75_138 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c139
+ bl_int_76_139 bl_int_75_139 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c140
+ bl_int_76_140 bl_int_75_140 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c141
+ bl_int_76_141 bl_int_75_141 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c142
+ bl_int_76_142 bl_int_75_142 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c143
+ bl_int_76_143 bl_int_75_143 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c144
+ bl_int_76_144 bl_int_75_144 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c145
+ bl_int_76_145 bl_int_75_145 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c146
+ bl_int_76_146 bl_int_75_146 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c147
+ bl_int_76_147 bl_int_75_147 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c148
+ bl_int_76_148 bl_int_75_148 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c149
+ bl_int_76_149 bl_int_75_149 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c150
+ bl_int_76_150 bl_int_75_150 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c151
+ bl_int_76_151 bl_int_75_151 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c152
+ bl_int_76_152 bl_int_75_152 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c153
+ bl_int_76_153 bl_int_75_153 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c154
+ bl_int_76_154 bl_int_75_154 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c155
+ bl_int_76_155 bl_int_75_155 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c156
+ bl_int_76_156 bl_int_75_156 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c157
+ bl_int_76_157 bl_int_75_157 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c158
+ bl_int_76_158 bl_int_75_158 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c159
+ bl_int_76_159 bl_int_75_159 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c160
+ bl_int_76_160 bl_int_75_160 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c161
+ bl_int_76_161 bl_int_75_161 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c162
+ bl_int_76_162 bl_int_75_162 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c163
+ bl_int_76_163 bl_int_75_163 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c164
+ bl_int_76_164 bl_int_75_164 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c165
+ bl_int_76_165 bl_int_75_165 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c166
+ bl_int_76_166 bl_int_75_166 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c167
+ bl_int_76_167 bl_int_75_167 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c168
+ bl_int_76_168 bl_int_75_168 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c169
+ bl_int_76_169 bl_int_75_169 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c170
+ bl_int_76_170 bl_int_75_170 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c171
+ bl_int_76_171 bl_int_75_171 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c172
+ bl_int_76_172 bl_int_75_172 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c173
+ bl_int_76_173 bl_int_75_173 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c174
+ bl_int_76_174 bl_int_75_174 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c175
+ bl_int_76_175 bl_int_75_175 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c176
+ bl_int_76_176 bl_int_75_176 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c177
+ bl_int_76_177 bl_int_75_177 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c178
+ bl_int_76_178 bl_int_75_178 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c179
+ bl_int_76_179 bl_int_75_179 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c180
+ bl_int_76_180 bl_int_75_180 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c181
+ bl_int_76_181 bl_int_75_181 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c182
+ bl_int_76_182 bl_int_75_182 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r76_c183
+ bl_int_76_183 bl_int_75_183 wl_0_76 gnd
+ sram_rom_base_one_cell
Xbit_r77_c0
+ bl_int_77_0 bl_int_76_0 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c1
+ bl_int_77_1 bl_int_76_1 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c2
+ bl_int_77_2 bl_int_76_2 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c3
+ bl_int_77_3 bl_int_76_3 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c4
+ bl_int_77_4 bl_int_76_4 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c5
+ bl_int_77_5 bl_int_76_5 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c6
+ bl_int_77_6 bl_int_76_6 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c7
+ bl_int_77_7 bl_int_76_7 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c8
+ bl_int_77_8 bl_int_76_8 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c9
+ bl_int_77_9 bl_int_76_9 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c10
+ bl_int_77_10 bl_int_76_10 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c11
+ bl_int_77_11 bl_int_76_11 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c12
+ bl_int_77_12 bl_int_76_12 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c13
+ bl_int_77_13 bl_int_76_13 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c14
+ bl_int_77_14 bl_int_76_14 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c15
+ bl_int_77_15 bl_int_76_15 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c16
+ bl_int_77_16 bl_int_76_16 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c17
+ bl_int_77_17 bl_int_76_17 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c18
+ bl_int_77_18 bl_int_76_18 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c19
+ bl_int_77_19 bl_int_76_19 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c20
+ bl_int_77_20 bl_int_76_20 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c21
+ bl_int_77_21 bl_int_76_21 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c22
+ bl_int_77_22 bl_int_76_22 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c23
+ bl_int_77_23 bl_int_76_23 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c24
+ bl_int_77_24 bl_int_76_24 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c25
+ bl_int_77_25 bl_int_76_25 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c26
+ bl_int_77_26 bl_int_76_26 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c27
+ bl_int_77_27 bl_int_76_27 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c28
+ bl_int_77_28 bl_int_76_28 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c29
+ bl_int_77_29 bl_int_76_29 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c30
+ bl_int_77_30 bl_int_76_30 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c31
+ bl_int_77_31 bl_int_76_31 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c32
+ bl_int_77_32 bl_int_76_32 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c33
+ bl_int_77_33 bl_int_76_33 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c34
+ bl_int_77_34 bl_int_76_34 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c35
+ bl_int_77_35 bl_int_76_35 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c36
+ bl_int_77_36 bl_int_76_36 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c37
+ bl_int_77_37 bl_int_76_37 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c38
+ bl_int_77_38 bl_int_76_38 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c39
+ bl_int_77_39 bl_int_76_39 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c40
+ bl_int_77_40 bl_int_76_40 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c41
+ bl_int_77_41 bl_int_76_41 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c42
+ bl_int_77_42 bl_int_76_42 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c43
+ bl_int_77_43 bl_int_76_43 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c44
+ bl_int_77_44 bl_int_76_44 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c45
+ bl_int_77_45 bl_int_76_45 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c46
+ bl_int_77_46 bl_int_76_46 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c47
+ bl_int_77_47 bl_int_76_47 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c48
+ bl_int_77_48 bl_int_76_48 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c49
+ bl_int_77_49 bl_int_76_49 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c50
+ bl_int_77_50 bl_int_76_50 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c51
+ bl_int_77_51 bl_int_76_51 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c52
+ bl_int_77_52 bl_int_76_52 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c53
+ bl_int_77_53 bl_int_76_53 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c54
+ bl_int_77_54 bl_int_76_54 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c55
+ bl_int_77_55 bl_int_76_55 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c56
+ bl_int_77_56 bl_int_76_56 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c57
+ bl_int_77_57 bl_int_76_57 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c58
+ bl_int_77_58 bl_int_76_58 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c59
+ bl_int_77_59 bl_int_76_59 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c60
+ bl_int_77_60 bl_int_76_60 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c61
+ bl_int_77_61 bl_int_76_61 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c62
+ bl_int_77_62 bl_int_76_62 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c63
+ bl_int_77_63 bl_int_76_63 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c64
+ bl_int_77_64 bl_int_76_64 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c65
+ bl_int_77_65 bl_int_76_65 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c66
+ bl_int_77_66 bl_int_76_66 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c67
+ bl_int_77_67 bl_int_76_67 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c68
+ bl_int_77_68 bl_int_76_68 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c69
+ bl_int_77_69 bl_int_76_69 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c70
+ bl_int_77_70 bl_int_76_70 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c71
+ bl_int_77_71 bl_int_76_71 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c72
+ bl_int_77_72 bl_int_76_72 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c73
+ bl_int_77_73 bl_int_76_73 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c74
+ bl_int_77_74 bl_int_76_74 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c75
+ bl_int_77_75 bl_int_76_75 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c76
+ bl_int_77_76 bl_int_76_76 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c77
+ bl_int_77_77 bl_int_76_77 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c78
+ bl_int_77_78 bl_int_76_78 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c79
+ bl_int_77_79 bl_int_76_79 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c80
+ bl_int_77_80 bl_int_76_80 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c81
+ bl_int_77_81 bl_int_76_81 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c82
+ bl_int_77_82 bl_int_76_82 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c83
+ bl_int_77_83 bl_int_76_83 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c84
+ bl_int_77_84 bl_int_76_84 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c85
+ bl_int_77_85 bl_int_76_85 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c86
+ bl_int_77_86 bl_int_76_86 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c87
+ bl_int_77_87 bl_int_76_87 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c88
+ bl_int_77_88 bl_int_76_88 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c89
+ bl_int_77_89 bl_int_76_89 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c90
+ bl_int_77_90 bl_int_76_90 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c91
+ bl_int_77_91 bl_int_76_91 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c92
+ bl_int_77_92 bl_int_76_92 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c93
+ bl_int_77_93 bl_int_76_93 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c94
+ bl_int_77_94 bl_int_76_94 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c95
+ bl_int_77_95 bl_int_76_95 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c96
+ bl_int_77_96 bl_int_76_96 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c97
+ bl_int_77_97 bl_int_76_97 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c98
+ bl_int_77_98 bl_int_76_98 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c99
+ bl_int_77_99 bl_int_76_99 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c100
+ bl_int_77_100 bl_int_76_100 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c101
+ bl_int_77_101 bl_int_76_101 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c102
+ bl_int_77_102 bl_int_76_102 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c103
+ bl_int_77_103 bl_int_76_103 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c104
+ bl_int_77_104 bl_int_76_104 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c105
+ bl_int_77_105 bl_int_76_105 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c106
+ bl_int_77_106 bl_int_76_106 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c107
+ bl_int_77_107 bl_int_76_107 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c108
+ bl_int_77_108 bl_int_76_108 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c109
+ bl_int_77_109 bl_int_76_109 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c110
+ bl_int_77_110 bl_int_76_110 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c111
+ bl_int_77_111 bl_int_76_111 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c112
+ bl_int_77_112 bl_int_76_112 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c113
+ bl_int_77_113 bl_int_76_113 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c114
+ bl_int_77_114 bl_int_76_114 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c115
+ bl_int_77_115 bl_int_76_115 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c116
+ bl_int_77_116 bl_int_76_116 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c117
+ bl_int_77_117 bl_int_76_117 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c118
+ bl_int_77_118 bl_int_76_118 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c119
+ bl_int_77_119 bl_int_76_119 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c120
+ bl_int_77_120 bl_int_76_120 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c121
+ bl_int_77_121 bl_int_76_121 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c122
+ bl_int_77_122 bl_int_76_122 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c123
+ bl_int_77_123 bl_int_76_123 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c124
+ bl_int_77_124 bl_int_76_124 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c125
+ bl_int_77_125 bl_int_76_125 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c126
+ bl_int_77_126 bl_int_76_126 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c127
+ bl_int_77_127 bl_int_76_127 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c128
+ bl_int_77_128 bl_int_76_128 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c129
+ bl_int_77_129 bl_int_76_129 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c130
+ bl_int_77_130 bl_int_76_130 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c131
+ bl_int_77_131 bl_int_76_131 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c132
+ bl_int_77_132 bl_int_76_132 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c133
+ bl_int_77_133 bl_int_76_133 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c134
+ bl_int_77_134 bl_int_76_134 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c135
+ bl_int_77_135 bl_int_76_135 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c136
+ bl_int_77_136 bl_int_76_136 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c137
+ bl_int_77_137 bl_int_76_137 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c138
+ bl_int_77_138 bl_int_76_138 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c139
+ bl_int_77_139 bl_int_76_139 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c140
+ bl_int_77_140 bl_int_76_140 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c141
+ bl_int_77_141 bl_int_76_141 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c142
+ bl_int_77_142 bl_int_76_142 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c143
+ bl_int_77_143 bl_int_76_143 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c144
+ bl_int_77_144 bl_int_76_144 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c145
+ bl_int_77_145 bl_int_76_145 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c146
+ bl_int_77_146 bl_int_76_146 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c147
+ bl_int_77_147 bl_int_76_147 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c148
+ bl_int_77_148 bl_int_76_148 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c149
+ bl_int_77_149 bl_int_76_149 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c150
+ bl_int_77_150 bl_int_76_150 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c151
+ bl_int_77_151 bl_int_76_151 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c152
+ bl_int_77_152 bl_int_76_152 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c153
+ bl_int_77_153 bl_int_76_153 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c154
+ bl_int_77_154 bl_int_76_154 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c155
+ bl_int_77_155 bl_int_76_155 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c156
+ bl_int_77_156 bl_int_76_156 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c157
+ bl_int_77_157 bl_int_76_157 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c158
+ bl_int_77_158 bl_int_76_158 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c159
+ bl_int_77_159 bl_int_76_159 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c160
+ bl_int_77_160 bl_int_76_160 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c161
+ bl_int_77_161 bl_int_76_161 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c162
+ bl_int_77_162 bl_int_76_162 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c163
+ bl_int_77_163 bl_int_76_163 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c164
+ bl_int_77_164 bl_int_76_164 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c165
+ bl_int_77_165 bl_int_76_165 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c166
+ bl_int_77_166 bl_int_76_166 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c167
+ bl_int_77_167 bl_int_76_167 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c168
+ bl_int_77_168 bl_int_76_168 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c169
+ bl_int_77_169 bl_int_76_169 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c170
+ bl_int_77_170 bl_int_76_170 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c171
+ bl_int_77_171 bl_int_76_171 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c172
+ bl_int_77_172 bl_int_76_172 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c173
+ bl_int_77_173 bl_int_76_173 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c174
+ bl_int_77_174 bl_int_76_174 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c175
+ bl_int_77_175 bl_int_76_175 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c176
+ bl_int_77_176 bl_int_76_176 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c177
+ bl_int_77_177 bl_int_76_177 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c178
+ bl_int_77_178 bl_int_76_178 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c179
+ bl_int_77_179 bl_int_76_179 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c180
+ bl_int_77_180 bl_int_76_180 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c181
+ bl_int_77_181 bl_int_76_181 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c182
+ bl_int_77_182 bl_int_76_182 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r77_c183
+ bl_int_77_183 bl_int_76_183 wl_0_77 gnd
+ sram_rom_base_one_cell
Xbit_r78_c0
+ bl_int_78_0 bl_int_77_0 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c1
+ bl_int_78_1 bl_int_77_1 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c2
+ bl_int_78_2 bl_int_77_2 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c3
+ bl_int_78_3 bl_int_77_3 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c4
+ bl_int_78_4 bl_int_77_4 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c5
+ bl_int_78_5 bl_int_77_5 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c6
+ bl_int_78_6 bl_int_77_6 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c7
+ bl_int_78_7 bl_int_77_7 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c8
+ bl_int_78_8 bl_int_77_8 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c9
+ bl_int_78_9 bl_int_77_9 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c10
+ bl_int_78_10 bl_int_77_10 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c11
+ bl_int_78_11 bl_int_77_11 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c12
+ bl_int_78_12 bl_int_77_12 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c13
+ bl_int_78_13 bl_int_77_13 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c14
+ bl_int_78_14 bl_int_77_14 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c15
+ bl_int_78_15 bl_int_77_15 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c16
+ bl_int_78_16 bl_int_77_16 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c17
+ bl_int_78_17 bl_int_77_17 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c18
+ bl_int_78_18 bl_int_77_18 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c19
+ bl_int_78_19 bl_int_77_19 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c20
+ bl_int_78_20 bl_int_77_20 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c21
+ bl_int_78_21 bl_int_77_21 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c22
+ bl_int_78_22 bl_int_77_22 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c23
+ bl_int_78_23 bl_int_77_23 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c24
+ bl_int_78_24 bl_int_77_24 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c25
+ bl_int_78_25 bl_int_77_25 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c26
+ bl_int_78_26 bl_int_77_26 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c27
+ bl_int_78_27 bl_int_77_27 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c28
+ bl_int_78_28 bl_int_77_28 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c29
+ bl_int_78_29 bl_int_77_29 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c30
+ bl_int_78_30 bl_int_77_30 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c31
+ bl_int_78_31 bl_int_77_31 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c32
+ bl_int_78_32 bl_int_77_32 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c33
+ bl_int_78_33 bl_int_77_33 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c34
+ bl_int_78_34 bl_int_77_34 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c35
+ bl_int_78_35 bl_int_77_35 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c36
+ bl_int_78_36 bl_int_77_36 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c37
+ bl_int_78_37 bl_int_77_37 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c38
+ bl_int_78_38 bl_int_77_38 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c39
+ bl_int_78_39 bl_int_77_39 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c40
+ bl_int_78_40 bl_int_77_40 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c41
+ bl_int_78_41 bl_int_77_41 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c42
+ bl_int_78_42 bl_int_77_42 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c43
+ bl_int_78_43 bl_int_77_43 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c44
+ bl_int_78_44 bl_int_77_44 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c45
+ bl_int_78_45 bl_int_77_45 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c46
+ bl_int_78_46 bl_int_77_46 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c47
+ bl_int_78_47 bl_int_77_47 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c48
+ bl_int_78_48 bl_int_77_48 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c49
+ bl_int_78_49 bl_int_77_49 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c50
+ bl_int_78_50 bl_int_77_50 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c51
+ bl_int_78_51 bl_int_77_51 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c52
+ bl_int_78_52 bl_int_77_52 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c53
+ bl_int_78_53 bl_int_77_53 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c54
+ bl_int_78_54 bl_int_77_54 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c55
+ bl_int_78_55 bl_int_77_55 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c56
+ bl_int_78_56 bl_int_77_56 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c57
+ bl_int_78_57 bl_int_77_57 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c58
+ bl_int_78_58 bl_int_77_58 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c59
+ bl_int_78_59 bl_int_77_59 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c60
+ bl_int_78_60 bl_int_77_60 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c61
+ bl_int_78_61 bl_int_77_61 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c62
+ bl_int_78_62 bl_int_77_62 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c63
+ bl_int_78_63 bl_int_77_63 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c64
+ bl_int_78_64 bl_int_77_64 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c65
+ bl_int_78_65 bl_int_77_65 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c66
+ bl_int_78_66 bl_int_77_66 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c67
+ bl_int_78_67 bl_int_77_67 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c68
+ bl_int_78_68 bl_int_77_68 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c69
+ bl_int_78_69 bl_int_77_69 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c70
+ bl_int_78_70 bl_int_77_70 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c71
+ bl_int_78_71 bl_int_77_71 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c72
+ bl_int_78_72 bl_int_77_72 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c73
+ bl_int_78_73 bl_int_77_73 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c74
+ bl_int_78_74 bl_int_77_74 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c75
+ bl_int_78_75 bl_int_77_75 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c76
+ bl_int_78_76 bl_int_77_76 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c77
+ bl_int_78_77 bl_int_77_77 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c78
+ bl_int_78_78 bl_int_77_78 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c79
+ bl_int_78_79 bl_int_77_79 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c80
+ bl_int_78_80 bl_int_77_80 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c81
+ bl_int_78_81 bl_int_77_81 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c82
+ bl_int_78_82 bl_int_77_82 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c83
+ bl_int_78_83 bl_int_77_83 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c84
+ bl_int_78_84 bl_int_77_84 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c85
+ bl_int_78_85 bl_int_77_85 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c86
+ bl_int_78_86 bl_int_77_86 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c87
+ bl_int_78_87 bl_int_77_87 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c88
+ bl_int_78_88 bl_int_77_88 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c89
+ bl_int_78_89 bl_int_77_89 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c90
+ bl_int_78_90 bl_int_77_90 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c91
+ bl_int_78_91 bl_int_77_91 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c92
+ bl_int_78_92 bl_int_77_92 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c93
+ bl_int_78_93 bl_int_77_93 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c94
+ bl_int_78_94 bl_int_77_94 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c95
+ bl_int_78_95 bl_int_77_95 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c96
+ bl_int_78_96 bl_int_77_96 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c97
+ bl_int_78_97 bl_int_77_97 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c98
+ bl_int_78_98 bl_int_77_98 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c99
+ bl_int_78_99 bl_int_77_99 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c100
+ bl_int_78_100 bl_int_77_100 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c101
+ bl_int_78_101 bl_int_77_101 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c102
+ bl_int_78_102 bl_int_77_102 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c103
+ bl_int_78_103 bl_int_77_103 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c104
+ bl_int_78_104 bl_int_77_104 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c105
+ bl_int_78_105 bl_int_77_105 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c106
+ bl_int_78_106 bl_int_77_106 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c107
+ bl_int_78_107 bl_int_77_107 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c108
+ bl_int_78_108 bl_int_77_108 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c109
+ bl_int_78_109 bl_int_77_109 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c110
+ bl_int_78_110 bl_int_77_110 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c111
+ bl_int_78_111 bl_int_77_111 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c112
+ bl_int_78_112 bl_int_77_112 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c113
+ bl_int_78_113 bl_int_77_113 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c114
+ bl_int_78_114 bl_int_77_114 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c115
+ bl_int_78_115 bl_int_77_115 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c116
+ bl_int_78_116 bl_int_77_116 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c117
+ bl_int_78_117 bl_int_77_117 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c118
+ bl_int_78_118 bl_int_77_118 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c119
+ bl_int_78_119 bl_int_77_119 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c120
+ bl_int_78_120 bl_int_77_120 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c121
+ bl_int_78_121 bl_int_77_121 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c122
+ bl_int_78_122 bl_int_77_122 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c123
+ bl_int_78_123 bl_int_77_123 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c124
+ bl_int_78_124 bl_int_77_124 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c125
+ bl_int_78_125 bl_int_77_125 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c126
+ bl_int_78_126 bl_int_77_126 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c127
+ bl_int_78_127 bl_int_77_127 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c128
+ bl_int_78_128 bl_int_77_128 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c129
+ bl_int_78_129 bl_int_77_129 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c130
+ bl_int_78_130 bl_int_77_130 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c131
+ bl_int_78_131 bl_int_77_131 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c132
+ bl_int_78_132 bl_int_77_132 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c133
+ bl_int_78_133 bl_int_77_133 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c134
+ bl_int_78_134 bl_int_77_134 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c135
+ bl_int_78_135 bl_int_77_135 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c136
+ bl_int_78_136 bl_int_77_136 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c137
+ bl_int_78_137 bl_int_77_137 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c138
+ bl_int_78_138 bl_int_77_138 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c139
+ bl_int_78_139 bl_int_77_139 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c140
+ bl_int_78_140 bl_int_77_140 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c141
+ bl_int_78_141 bl_int_77_141 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c142
+ bl_int_78_142 bl_int_77_142 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c143
+ bl_int_78_143 bl_int_77_143 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c144
+ bl_int_78_144 bl_int_77_144 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c145
+ bl_int_78_145 bl_int_77_145 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c146
+ bl_int_78_146 bl_int_77_146 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c147
+ bl_int_78_147 bl_int_77_147 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c148
+ bl_int_78_148 bl_int_77_148 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c149
+ bl_int_78_149 bl_int_77_149 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c150
+ bl_int_78_150 bl_int_77_150 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c151
+ bl_int_78_151 bl_int_77_151 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c152
+ bl_int_78_152 bl_int_77_152 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c153
+ bl_int_78_153 bl_int_77_153 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c154
+ bl_int_78_154 bl_int_77_154 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c155
+ bl_int_78_155 bl_int_77_155 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c156
+ bl_int_78_156 bl_int_77_156 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c157
+ bl_int_78_157 bl_int_77_157 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c158
+ bl_int_78_158 bl_int_77_158 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c159
+ bl_int_78_159 bl_int_77_159 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c160
+ bl_int_78_160 bl_int_77_160 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c161
+ bl_int_78_161 bl_int_77_161 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c162
+ bl_int_78_162 bl_int_77_162 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c163
+ bl_int_78_163 bl_int_77_163 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c164
+ bl_int_78_164 bl_int_77_164 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c165
+ bl_int_78_165 bl_int_77_165 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c166
+ bl_int_78_166 bl_int_77_166 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c167
+ bl_int_78_167 bl_int_77_167 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c168
+ bl_int_78_168 bl_int_77_168 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c169
+ bl_int_78_169 bl_int_77_169 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c170
+ bl_int_78_170 bl_int_77_170 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c171
+ bl_int_78_171 bl_int_77_171 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c172
+ bl_int_78_172 bl_int_77_172 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c173
+ bl_int_78_173 bl_int_77_173 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c174
+ bl_int_78_174 bl_int_77_174 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c175
+ bl_int_78_175 bl_int_77_175 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c176
+ bl_int_78_176 bl_int_77_176 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c177
+ bl_int_78_177 bl_int_77_177 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c178
+ bl_int_78_178 bl_int_77_178 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c179
+ bl_int_78_179 bl_int_77_179 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c180
+ bl_int_78_180 bl_int_77_180 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c181
+ bl_int_78_181 bl_int_77_181 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c182
+ bl_int_78_182 bl_int_77_182 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r78_c183
+ bl_int_78_183 bl_int_77_183 wl_0_78 gnd
+ sram_rom_base_one_cell
Xbit_r79_c0
+ bl_int_79_0 bl_int_78_0 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c1
+ bl_int_79_1 bl_int_78_1 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c2
+ bl_int_79_2 bl_int_78_2 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c3
+ bl_int_79_3 bl_int_78_3 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c4
+ bl_int_79_4 bl_int_78_4 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c5
+ bl_int_79_5 bl_int_78_5 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c6
+ bl_int_79_6 bl_int_78_6 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c7
+ bl_int_79_7 bl_int_78_7 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c8
+ bl_int_79_8 bl_int_78_8 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c9
+ bl_int_79_9 bl_int_78_9 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c10
+ bl_int_79_10 bl_int_78_10 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c11
+ bl_int_79_11 bl_int_78_11 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c12
+ bl_int_79_12 bl_int_78_12 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c13
+ bl_int_79_13 bl_int_78_13 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c14
+ bl_int_79_14 bl_int_78_14 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c15
+ bl_int_79_15 bl_int_78_15 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c16
+ bl_int_79_16 bl_int_78_16 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c17
+ bl_int_79_17 bl_int_78_17 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c18
+ bl_int_79_18 bl_int_78_18 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c19
+ bl_int_79_19 bl_int_78_19 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c20
+ bl_int_79_20 bl_int_78_20 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c21
+ bl_int_79_21 bl_int_78_21 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c22
+ bl_int_79_22 bl_int_78_22 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c23
+ bl_int_79_23 bl_int_78_23 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c24
+ bl_int_79_24 bl_int_78_24 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c25
+ bl_int_79_25 bl_int_78_25 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c26
+ bl_int_79_26 bl_int_78_26 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c27
+ bl_int_79_27 bl_int_78_27 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c28
+ bl_int_79_28 bl_int_78_28 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c29
+ bl_int_79_29 bl_int_78_29 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c30
+ bl_int_79_30 bl_int_78_30 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c31
+ bl_int_79_31 bl_int_78_31 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c32
+ bl_int_79_32 bl_int_78_32 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c33
+ bl_int_79_33 bl_int_78_33 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c34
+ bl_int_79_34 bl_int_78_34 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c35
+ bl_int_79_35 bl_int_78_35 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c36
+ bl_int_79_36 bl_int_78_36 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c37
+ bl_int_79_37 bl_int_78_37 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c38
+ bl_int_79_38 bl_int_78_38 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c39
+ bl_int_79_39 bl_int_78_39 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c40
+ bl_int_79_40 bl_int_78_40 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c41
+ bl_int_79_41 bl_int_78_41 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c42
+ bl_int_79_42 bl_int_78_42 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c43
+ bl_int_79_43 bl_int_78_43 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c44
+ bl_int_79_44 bl_int_78_44 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c45
+ bl_int_79_45 bl_int_78_45 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c46
+ bl_int_79_46 bl_int_78_46 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c47
+ bl_int_79_47 bl_int_78_47 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c48
+ bl_int_79_48 bl_int_78_48 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c49
+ bl_int_79_49 bl_int_78_49 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c50
+ bl_int_79_50 bl_int_78_50 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c51
+ bl_int_79_51 bl_int_78_51 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c52
+ bl_int_79_52 bl_int_78_52 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c53
+ bl_int_79_53 bl_int_78_53 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c54
+ bl_int_79_54 bl_int_78_54 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c55
+ bl_int_79_55 bl_int_78_55 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c56
+ bl_int_79_56 bl_int_78_56 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c57
+ bl_int_79_57 bl_int_78_57 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c58
+ bl_int_79_58 bl_int_78_58 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c59
+ bl_int_79_59 bl_int_78_59 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c60
+ bl_int_79_60 bl_int_78_60 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c61
+ bl_int_79_61 bl_int_78_61 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c62
+ bl_int_79_62 bl_int_78_62 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c63
+ bl_int_79_63 bl_int_78_63 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c64
+ bl_int_79_64 bl_int_78_64 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c65
+ bl_int_79_65 bl_int_78_65 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c66
+ bl_int_79_66 bl_int_78_66 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c67
+ bl_int_79_67 bl_int_78_67 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c68
+ bl_int_79_68 bl_int_78_68 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c69
+ bl_int_79_69 bl_int_78_69 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c70
+ bl_int_79_70 bl_int_78_70 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c71
+ bl_int_79_71 bl_int_78_71 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c72
+ bl_int_79_72 bl_int_78_72 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c73
+ bl_int_79_73 bl_int_78_73 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c74
+ bl_int_79_74 bl_int_78_74 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c75
+ bl_int_79_75 bl_int_78_75 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c76
+ bl_int_79_76 bl_int_78_76 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c77
+ bl_int_79_77 bl_int_78_77 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c78
+ bl_int_79_78 bl_int_78_78 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c79
+ bl_int_79_79 bl_int_78_79 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c80
+ bl_int_79_80 bl_int_78_80 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c81
+ bl_int_79_81 bl_int_78_81 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c82
+ bl_int_79_82 bl_int_78_82 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c83
+ bl_int_79_83 bl_int_78_83 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c84
+ bl_int_79_84 bl_int_78_84 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c85
+ bl_int_79_85 bl_int_78_85 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c86
+ bl_int_79_86 bl_int_78_86 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c87
+ bl_int_79_87 bl_int_78_87 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c88
+ bl_int_79_88 bl_int_78_88 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c89
+ bl_int_79_89 bl_int_78_89 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c90
+ bl_int_79_90 bl_int_78_90 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c91
+ bl_int_79_91 bl_int_78_91 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c92
+ bl_int_79_92 bl_int_78_92 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c93
+ bl_int_79_93 bl_int_78_93 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c94
+ bl_int_79_94 bl_int_78_94 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c95
+ bl_int_79_95 bl_int_78_95 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c96
+ bl_int_79_96 bl_int_78_96 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c97
+ bl_int_79_97 bl_int_78_97 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c98
+ bl_int_79_98 bl_int_78_98 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c99
+ bl_int_79_99 bl_int_78_99 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c100
+ bl_int_79_100 bl_int_78_100 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c101
+ bl_int_79_101 bl_int_78_101 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c102
+ bl_int_79_102 bl_int_78_102 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c103
+ bl_int_79_103 bl_int_78_103 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c104
+ bl_int_79_104 bl_int_78_104 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c105
+ bl_int_79_105 bl_int_78_105 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c106
+ bl_int_79_106 bl_int_78_106 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c107
+ bl_int_79_107 bl_int_78_107 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c108
+ bl_int_79_108 bl_int_78_108 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c109
+ bl_int_79_109 bl_int_78_109 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c110
+ bl_int_79_110 bl_int_78_110 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c111
+ bl_int_79_111 bl_int_78_111 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c112
+ bl_int_79_112 bl_int_78_112 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c113
+ bl_int_79_113 bl_int_78_113 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c114
+ bl_int_79_114 bl_int_78_114 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c115
+ bl_int_79_115 bl_int_78_115 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c116
+ bl_int_79_116 bl_int_78_116 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c117
+ bl_int_79_117 bl_int_78_117 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c118
+ bl_int_79_118 bl_int_78_118 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c119
+ bl_int_79_119 bl_int_78_119 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c120
+ bl_int_79_120 bl_int_78_120 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c121
+ bl_int_79_121 bl_int_78_121 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c122
+ bl_int_79_122 bl_int_78_122 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c123
+ bl_int_79_123 bl_int_78_123 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c124
+ bl_int_79_124 bl_int_78_124 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c125
+ bl_int_79_125 bl_int_78_125 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c126
+ bl_int_79_126 bl_int_78_126 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c127
+ bl_int_79_127 bl_int_78_127 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c128
+ bl_int_79_128 bl_int_78_128 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c129
+ bl_int_79_129 bl_int_78_129 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c130
+ bl_int_79_130 bl_int_78_130 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c131
+ bl_int_79_131 bl_int_78_131 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c132
+ bl_int_79_132 bl_int_78_132 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c133
+ bl_int_79_133 bl_int_78_133 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c134
+ bl_int_79_134 bl_int_78_134 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c135
+ bl_int_79_135 bl_int_78_135 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c136
+ bl_int_79_136 bl_int_78_136 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c137
+ bl_int_79_137 bl_int_78_137 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c138
+ bl_int_79_138 bl_int_78_138 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c139
+ bl_int_79_139 bl_int_78_139 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c140
+ bl_int_79_140 bl_int_78_140 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c141
+ bl_int_79_141 bl_int_78_141 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c142
+ bl_int_79_142 bl_int_78_142 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c143
+ bl_int_79_143 bl_int_78_143 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c144
+ bl_int_79_144 bl_int_78_144 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c145
+ bl_int_79_145 bl_int_78_145 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c146
+ bl_int_79_146 bl_int_78_146 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c147
+ bl_int_79_147 bl_int_78_147 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c148
+ bl_int_79_148 bl_int_78_148 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c149
+ bl_int_79_149 bl_int_78_149 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c150
+ bl_int_79_150 bl_int_78_150 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c151
+ bl_int_79_151 bl_int_78_151 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c152
+ bl_int_79_152 bl_int_78_152 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c153
+ bl_int_79_153 bl_int_78_153 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c154
+ bl_int_79_154 bl_int_78_154 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c155
+ bl_int_79_155 bl_int_78_155 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c156
+ bl_int_79_156 bl_int_78_156 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c157
+ bl_int_79_157 bl_int_78_157 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c158
+ bl_int_79_158 bl_int_78_158 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c159
+ bl_int_79_159 bl_int_78_159 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c160
+ bl_int_79_160 bl_int_78_160 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c161
+ bl_int_79_161 bl_int_78_161 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c162
+ bl_int_79_162 bl_int_78_162 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c163
+ bl_int_79_163 bl_int_78_163 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c164
+ bl_int_79_164 bl_int_78_164 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c165
+ bl_int_79_165 bl_int_78_165 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c166
+ bl_int_79_166 bl_int_78_166 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c167
+ bl_int_79_167 bl_int_78_167 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c168
+ bl_int_79_168 bl_int_78_168 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c169
+ bl_int_79_169 bl_int_78_169 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c170
+ bl_int_79_170 bl_int_78_170 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c171
+ bl_int_79_171 bl_int_78_171 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c172
+ bl_int_79_172 bl_int_78_172 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c173
+ bl_int_79_173 bl_int_78_173 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c174
+ bl_int_79_174 bl_int_78_174 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c175
+ bl_int_79_175 bl_int_78_175 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c176
+ bl_int_79_176 bl_int_78_176 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c177
+ bl_int_79_177 bl_int_78_177 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c178
+ bl_int_79_178 bl_int_78_178 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c179
+ bl_int_79_179 bl_int_78_179 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c180
+ bl_int_79_180 bl_int_78_180 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c181
+ bl_int_79_181 bl_int_78_181 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c182
+ bl_int_79_182 bl_int_78_182 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r79_c183
+ bl_int_79_183 bl_int_78_183 wl_0_79 gnd
+ sram_rom_base_one_cell
Xbit_r80_c0
+ bl_int_80_0 bl_int_79_0 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c1
+ bl_int_80_1 bl_int_79_1 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c2
+ bl_int_80_2 bl_int_79_2 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c3
+ bl_int_80_3 bl_int_79_3 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c4
+ bl_int_80_4 bl_int_79_4 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c5
+ bl_int_80_5 bl_int_79_5 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c6
+ bl_int_80_6 bl_int_79_6 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c7
+ bl_int_80_7 bl_int_79_7 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c8
+ bl_int_80_8 bl_int_79_8 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c9
+ bl_int_80_9 bl_int_79_9 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c10
+ bl_int_80_10 bl_int_79_10 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c11
+ bl_int_80_11 bl_int_79_11 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c12
+ bl_int_80_12 bl_int_79_12 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c13
+ bl_int_80_13 bl_int_79_13 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c14
+ bl_int_80_14 bl_int_79_14 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c15
+ bl_int_80_15 bl_int_79_15 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c16
+ bl_int_80_16 bl_int_79_16 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c17
+ bl_int_80_17 bl_int_79_17 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c18
+ bl_int_80_18 bl_int_79_18 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c19
+ bl_int_80_19 bl_int_79_19 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c20
+ bl_int_80_20 bl_int_79_20 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c21
+ bl_int_80_21 bl_int_79_21 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c22
+ bl_int_80_22 bl_int_79_22 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c23
+ bl_int_80_23 bl_int_79_23 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c24
+ bl_int_80_24 bl_int_79_24 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c25
+ bl_int_80_25 bl_int_79_25 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c26
+ bl_int_80_26 bl_int_79_26 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c27
+ bl_int_80_27 bl_int_79_27 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c28
+ bl_int_80_28 bl_int_79_28 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c29
+ bl_int_80_29 bl_int_79_29 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c30
+ bl_int_80_30 bl_int_79_30 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c31
+ bl_int_80_31 bl_int_79_31 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c32
+ bl_int_80_32 bl_int_79_32 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c33
+ bl_int_80_33 bl_int_79_33 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c34
+ bl_int_80_34 bl_int_79_34 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c35
+ bl_int_80_35 bl_int_79_35 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c36
+ bl_int_80_36 bl_int_79_36 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c37
+ bl_int_80_37 bl_int_79_37 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c38
+ bl_int_80_38 bl_int_79_38 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c39
+ bl_int_80_39 bl_int_79_39 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c40
+ bl_int_80_40 bl_int_79_40 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c41
+ bl_int_80_41 bl_int_79_41 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c42
+ bl_int_80_42 bl_int_79_42 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c43
+ bl_int_80_43 bl_int_79_43 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c44
+ bl_int_80_44 bl_int_79_44 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c45
+ bl_int_80_45 bl_int_79_45 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c46
+ bl_int_80_46 bl_int_79_46 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c47
+ bl_int_80_47 bl_int_79_47 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c48
+ bl_int_80_48 bl_int_79_48 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c49
+ bl_int_80_49 bl_int_79_49 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c50
+ bl_int_80_50 bl_int_79_50 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c51
+ bl_int_80_51 bl_int_79_51 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c52
+ bl_int_80_52 bl_int_79_52 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c53
+ bl_int_80_53 bl_int_79_53 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c54
+ bl_int_80_54 bl_int_79_54 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c55
+ bl_int_80_55 bl_int_79_55 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c56
+ bl_int_80_56 bl_int_79_56 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c57
+ bl_int_80_57 bl_int_79_57 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c58
+ bl_int_80_58 bl_int_79_58 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c59
+ bl_int_80_59 bl_int_79_59 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c60
+ bl_int_80_60 bl_int_79_60 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c61
+ bl_int_80_61 bl_int_79_61 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c62
+ bl_int_80_62 bl_int_79_62 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c63
+ bl_int_80_63 bl_int_79_63 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c64
+ bl_int_80_64 bl_int_79_64 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c65
+ bl_int_80_65 bl_int_79_65 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c66
+ bl_int_80_66 bl_int_79_66 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c67
+ bl_int_80_67 bl_int_79_67 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c68
+ bl_int_80_68 bl_int_79_68 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c69
+ bl_int_80_69 bl_int_79_69 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c70
+ bl_int_80_70 bl_int_79_70 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c71
+ bl_int_80_71 bl_int_79_71 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c72
+ bl_int_80_72 bl_int_79_72 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c73
+ bl_int_80_73 bl_int_79_73 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c74
+ bl_int_80_74 bl_int_79_74 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c75
+ bl_int_80_75 bl_int_79_75 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c76
+ bl_int_80_76 bl_int_79_76 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c77
+ bl_int_80_77 bl_int_79_77 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c78
+ bl_int_80_78 bl_int_79_78 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c79
+ bl_int_80_79 bl_int_79_79 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c80
+ bl_int_80_80 bl_int_79_80 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c81
+ bl_int_80_81 bl_int_79_81 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c82
+ bl_int_80_82 bl_int_79_82 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c83
+ bl_int_80_83 bl_int_79_83 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c84
+ bl_int_80_84 bl_int_79_84 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c85
+ bl_int_80_85 bl_int_79_85 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c86
+ bl_int_80_86 bl_int_79_86 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c87
+ bl_int_80_87 bl_int_79_87 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c88
+ bl_int_80_88 bl_int_79_88 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c89
+ bl_int_80_89 bl_int_79_89 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c90
+ bl_int_80_90 bl_int_79_90 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c91
+ bl_int_80_91 bl_int_79_91 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c92
+ bl_int_80_92 bl_int_79_92 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c93
+ bl_int_80_93 bl_int_79_93 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c94
+ bl_int_80_94 bl_int_79_94 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c95
+ bl_int_80_95 bl_int_79_95 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c96
+ bl_int_80_96 bl_int_79_96 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c97
+ bl_int_80_97 bl_int_79_97 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c98
+ bl_int_80_98 bl_int_79_98 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c99
+ bl_int_80_99 bl_int_79_99 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c100
+ bl_int_80_100 bl_int_79_100 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c101
+ bl_int_80_101 bl_int_79_101 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c102
+ bl_int_80_102 bl_int_79_102 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c103
+ bl_int_80_103 bl_int_79_103 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c104
+ bl_int_80_104 bl_int_79_104 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c105
+ bl_int_80_105 bl_int_79_105 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c106
+ bl_int_80_106 bl_int_79_106 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c107
+ bl_int_80_107 bl_int_79_107 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c108
+ bl_int_80_108 bl_int_79_108 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c109
+ bl_int_80_109 bl_int_79_109 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c110
+ bl_int_80_110 bl_int_79_110 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c111
+ bl_int_80_111 bl_int_79_111 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c112
+ bl_int_80_112 bl_int_79_112 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c113
+ bl_int_80_113 bl_int_79_113 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c114
+ bl_int_80_114 bl_int_79_114 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c115
+ bl_int_80_115 bl_int_79_115 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c116
+ bl_int_80_116 bl_int_79_116 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c117
+ bl_int_80_117 bl_int_79_117 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c118
+ bl_int_80_118 bl_int_79_118 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c119
+ bl_int_80_119 bl_int_79_119 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c120
+ bl_int_80_120 bl_int_79_120 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c121
+ bl_int_80_121 bl_int_79_121 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c122
+ bl_int_80_122 bl_int_79_122 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c123
+ bl_int_80_123 bl_int_79_123 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c124
+ bl_int_80_124 bl_int_79_124 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c125
+ bl_int_80_125 bl_int_79_125 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c126
+ bl_int_80_126 bl_int_79_126 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c127
+ bl_int_80_127 bl_int_79_127 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c128
+ bl_int_80_128 bl_int_79_128 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c129
+ bl_int_80_129 bl_int_79_129 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c130
+ bl_int_80_130 bl_int_79_130 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c131
+ bl_int_80_131 bl_int_79_131 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c132
+ bl_int_80_132 bl_int_79_132 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c133
+ bl_int_80_133 bl_int_79_133 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c134
+ bl_int_80_134 bl_int_79_134 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c135
+ bl_int_80_135 bl_int_79_135 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c136
+ bl_int_80_136 bl_int_79_136 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c137
+ bl_int_80_137 bl_int_79_137 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c138
+ bl_int_80_138 bl_int_79_138 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c139
+ bl_int_80_139 bl_int_79_139 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c140
+ bl_int_80_140 bl_int_79_140 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c141
+ bl_int_80_141 bl_int_79_141 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c142
+ bl_int_80_142 bl_int_79_142 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c143
+ bl_int_80_143 bl_int_79_143 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c144
+ bl_int_80_144 bl_int_79_144 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c145
+ bl_int_80_145 bl_int_79_145 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c146
+ bl_int_80_146 bl_int_79_146 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c147
+ bl_int_80_147 bl_int_79_147 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c148
+ bl_int_80_148 bl_int_79_148 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c149
+ bl_int_80_149 bl_int_79_149 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c150
+ bl_int_80_150 bl_int_79_150 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c151
+ bl_int_80_151 bl_int_79_151 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c152
+ bl_int_80_152 bl_int_79_152 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c153
+ bl_int_80_153 bl_int_79_153 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c154
+ bl_int_80_154 bl_int_79_154 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c155
+ bl_int_80_155 bl_int_79_155 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c156
+ bl_int_80_156 bl_int_79_156 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c157
+ bl_int_80_157 bl_int_79_157 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c158
+ bl_int_80_158 bl_int_79_158 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c159
+ bl_int_80_159 bl_int_79_159 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c160
+ bl_int_80_160 bl_int_79_160 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c161
+ bl_int_80_161 bl_int_79_161 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c162
+ bl_int_80_162 bl_int_79_162 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c163
+ bl_int_80_163 bl_int_79_163 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c164
+ bl_int_80_164 bl_int_79_164 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c165
+ bl_int_80_165 bl_int_79_165 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c166
+ bl_int_80_166 bl_int_79_166 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c167
+ bl_int_80_167 bl_int_79_167 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c168
+ bl_int_80_168 bl_int_79_168 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c169
+ bl_int_80_169 bl_int_79_169 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c170
+ bl_int_80_170 bl_int_79_170 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c171
+ bl_int_80_171 bl_int_79_171 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c172
+ bl_int_80_172 bl_int_79_172 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c173
+ bl_int_80_173 bl_int_79_173 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c174
+ bl_int_80_174 bl_int_79_174 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c175
+ bl_int_80_175 bl_int_79_175 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c176
+ bl_int_80_176 bl_int_79_176 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c177
+ bl_int_80_177 bl_int_79_177 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c178
+ bl_int_80_178 bl_int_79_178 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c179
+ bl_int_80_179 bl_int_79_179 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c180
+ bl_int_80_180 bl_int_79_180 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c181
+ bl_int_80_181 bl_int_79_181 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c182
+ bl_int_80_182 bl_int_79_182 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r80_c183
+ bl_int_80_183 bl_int_79_183 wl_0_80 gnd
+ sram_rom_base_one_cell
Xbit_r81_c0
+ bl_int_81_0 bl_int_80_0 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c1
+ bl_int_81_1 bl_int_80_1 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c2
+ bl_int_81_2 bl_int_80_2 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c3
+ bl_int_81_3 bl_int_80_3 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c4
+ bl_int_81_4 bl_int_80_4 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c5
+ bl_int_81_5 bl_int_80_5 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c6
+ bl_int_81_6 bl_int_80_6 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c7
+ bl_int_81_7 bl_int_80_7 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c8
+ bl_int_81_8 bl_int_80_8 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c9
+ bl_int_81_9 bl_int_80_9 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c10
+ bl_int_81_10 bl_int_80_10 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c11
+ bl_int_81_11 bl_int_80_11 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c12
+ bl_int_81_12 bl_int_80_12 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c13
+ bl_int_81_13 bl_int_80_13 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c14
+ bl_int_81_14 bl_int_80_14 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c15
+ bl_int_81_15 bl_int_80_15 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c16
+ bl_int_81_16 bl_int_80_16 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c17
+ bl_int_81_17 bl_int_80_17 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c18
+ bl_int_81_18 bl_int_80_18 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c19
+ bl_int_81_19 bl_int_80_19 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c20
+ bl_int_81_20 bl_int_80_20 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c21
+ bl_int_81_21 bl_int_80_21 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c22
+ bl_int_81_22 bl_int_80_22 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c23
+ bl_int_81_23 bl_int_80_23 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c24
+ bl_int_81_24 bl_int_80_24 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c25
+ bl_int_81_25 bl_int_80_25 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c26
+ bl_int_81_26 bl_int_80_26 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c27
+ bl_int_81_27 bl_int_80_27 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c28
+ bl_int_81_28 bl_int_80_28 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c29
+ bl_int_81_29 bl_int_80_29 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c30
+ bl_int_81_30 bl_int_80_30 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c31
+ bl_int_81_31 bl_int_80_31 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c32
+ bl_int_81_32 bl_int_80_32 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c33
+ bl_int_81_33 bl_int_80_33 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c34
+ bl_int_81_34 bl_int_80_34 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c35
+ bl_int_81_35 bl_int_80_35 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c36
+ bl_int_81_36 bl_int_80_36 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c37
+ bl_int_81_37 bl_int_80_37 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c38
+ bl_int_81_38 bl_int_80_38 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c39
+ bl_int_81_39 bl_int_80_39 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c40
+ bl_int_81_40 bl_int_80_40 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c41
+ bl_int_81_41 bl_int_80_41 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c42
+ bl_int_81_42 bl_int_80_42 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c43
+ bl_int_81_43 bl_int_80_43 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c44
+ bl_int_81_44 bl_int_80_44 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c45
+ bl_int_81_45 bl_int_80_45 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c46
+ bl_int_81_46 bl_int_80_46 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c47
+ bl_int_81_47 bl_int_80_47 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c48
+ bl_int_81_48 bl_int_80_48 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c49
+ bl_int_81_49 bl_int_80_49 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c50
+ bl_int_81_50 bl_int_80_50 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c51
+ bl_int_81_51 bl_int_80_51 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c52
+ bl_int_81_52 bl_int_80_52 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c53
+ bl_int_81_53 bl_int_80_53 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c54
+ bl_int_81_54 bl_int_80_54 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c55
+ bl_int_81_55 bl_int_80_55 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c56
+ bl_int_81_56 bl_int_80_56 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c57
+ bl_int_81_57 bl_int_80_57 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c58
+ bl_int_81_58 bl_int_80_58 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c59
+ bl_int_81_59 bl_int_80_59 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c60
+ bl_int_81_60 bl_int_80_60 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c61
+ bl_int_81_61 bl_int_80_61 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c62
+ bl_int_81_62 bl_int_80_62 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c63
+ bl_int_81_63 bl_int_80_63 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c64
+ bl_int_81_64 bl_int_80_64 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c65
+ bl_int_81_65 bl_int_80_65 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c66
+ bl_int_81_66 bl_int_80_66 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c67
+ bl_int_81_67 bl_int_80_67 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c68
+ bl_int_81_68 bl_int_80_68 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c69
+ bl_int_81_69 bl_int_80_69 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c70
+ bl_int_81_70 bl_int_80_70 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c71
+ bl_int_81_71 bl_int_80_71 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c72
+ bl_int_81_72 bl_int_80_72 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c73
+ bl_int_81_73 bl_int_80_73 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c74
+ bl_int_81_74 bl_int_80_74 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c75
+ bl_int_81_75 bl_int_80_75 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c76
+ bl_int_81_76 bl_int_80_76 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c77
+ bl_int_81_77 bl_int_80_77 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c78
+ bl_int_81_78 bl_int_80_78 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c79
+ bl_int_81_79 bl_int_80_79 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c80
+ bl_int_81_80 bl_int_80_80 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c81
+ bl_int_81_81 bl_int_80_81 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c82
+ bl_int_81_82 bl_int_80_82 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c83
+ bl_int_81_83 bl_int_80_83 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c84
+ bl_int_81_84 bl_int_80_84 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c85
+ bl_int_81_85 bl_int_80_85 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c86
+ bl_int_81_86 bl_int_80_86 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c87
+ bl_int_81_87 bl_int_80_87 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c88
+ bl_int_81_88 bl_int_80_88 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c89
+ bl_int_81_89 bl_int_80_89 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c90
+ bl_int_81_90 bl_int_80_90 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c91
+ bl_int_81_91 bl_int_80_91 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c92
+ bl_int_81_92 bl_int_80_92 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c93
+ bl_int_81_93 bl_int_80_93 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c94
+ bl_int_81_94 bl_int_80_94 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c95
+ bl_int_81_95 bl_int_80_95 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c96
+ bl_int_81_96 bl_int_80_96 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c97
+ bl_int_81_97 bl_int_80_97 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c98
+ bl_int_81_98 bl_int_80_98 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c99
+ bl_int_81_99 bl_int_80_99 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c100
+ bl_int_81_100 bl_int_80_100 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c101
+ bl_int_81_101 bl_int_80_101 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c102
+ bl_int_81_102 bl_int_80_102 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c103
+ bl_int_81_103 bl_int_80_103 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c104
+ bl_int_81_104 bl_int_80_104 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c105
+ bl_int_81_105 bl_int_80_105 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c106
+ bl_int_81_106 bl_int_80_106 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c107
+ bl_int_81_107 bl_int_80_107 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c108
+ bl_int_81_108 bl_int_80_108 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c109
+ bl_int_81_109 bl_int_80_109 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c110
+ bl_int_81_110 bl_int_80_110 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c111
+ bl_int_81_111 bl_int_80_111 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c112
+ bl_int_81_112 bl_int_80_112 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c113
+ bl_int_81_113 bl_int_80_113 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c114
+ bl_int_81_114 bl_int_80_114 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c115
+ bl_int_81_115 bl_int_80_115 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c116
+ bl_int_81_116 bl_int_80_116 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c117
+ bl_int_81_117 bl_int_80_117 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c118
+ bl_int_81_118 bl_int_80_118 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c119
+ bl_int_81_119 bl_int_80_119 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c120
+ bl_int_81_120 bl_int_80_120 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c121
+ bl_int_81_121 bl_int_80_121 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c122
+ bl_int_81_122 bl_int_80_122 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c123
+ bl_int_81_123 bl_int_80_123 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c124
+ bl_int_81_124 bl_int_80_124 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c125
+ bl_int_81_125 bl_int_80_125 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c126
+ bl_int_81_126 bl_int_80_126 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c127
+ bl_int_81_127 bl_int_80_127 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c128
+ bl_int_81_128 bl_int_80_128 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c129
+ bl_int_81_129 bl_int_80_129 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c130
+ bl_int_81_130 bl_int_80_130 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c131
+ bl_int_81_131 bl_int_80_131 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c132
+ bl_int_81_132 bl_int_80_132 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c133
+ bl_int_81_133 bl_int_80_133 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c134
+ bl_int_81_134 bl_int_80_134 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c135
+ bl_int_81_135 bl_int_80_135 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c136
+ bl_int_81_136 bl_int_80_136 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c137
+ bl_int_81_137 bl_int_80_137 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c138
+ bl_int_81_138 bl_int_80_138 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c139
+ bl_int_81_139 bl_int_80_139 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c140
+ bl_int_81_140 bl_int_80_140 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c141
+ bl_int_81_141 bl_int_80_141 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c142
+ bl_int_81_142 bl_int_80_142 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c143
+ bl_int_81_143 bl_int_80_143 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c144
+ bl_int_81_144 bl_int_80_144 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c145
+ bl_int_81_145 bl_int_80_145 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c146
+ bl_int_81_146 bl_int_80_146 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c147
+ bl_int_81_147 bl_int_80_147 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c148
+ bl_int_81_148 bl_int_80_148 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c149
+ bl_int_81_149 bl_int_80_149 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c150
+ bl_int_81_150 bl_int_80_150 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c151
+ bl_int_81_151 bl_int_80_151 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c152
+ bl_int_81_152 bl_int_80_152 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c153
+ bl_int_81_153 bl_int_80_153 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c154
+ bl_int_81_154 bl_int_80_154 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c155
+ bl_int_81_155 bl_int_80_155 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c156
+ bl_int_81_156 bl_int_80_156 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c157
+ bl_int_81_157 bl_int_80_157 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c158
+ bl_int_81_158 bl_int_80_158 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c159
+ bl_int_81_159 bl_int_80_159 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c160
+ bl_int_81_160 bl_int_80_160 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c161
+ bl_int_81_161 bl_int_80_161 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c162
+ bl_int_81_162 bl_int_80_162 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c163
+ bl_int_81_163 bl_int_80_163 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c164
+ bl_int_81_164 bl_int_80_164 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c165
+ bl_int_81_165 bl_int_80_165 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c166
+ bl_int_81_166 bl_int_80_166 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c167
+ bl_int_81_167 bl_int_80_167 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c168
+ bl_int_81_168 bl_int_80_168 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c169
+ bl_int_81_169 bl_int_80_169 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c170
+ bl_int_81_170 bl_int_80_170 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c171
+ bl_int_81_171 bl_int_80_171 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c172
+ bl_int_81_172 bl_int_80_172 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c173
+ bl_int_81_173 bl_int_80_173 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c174
+ bl_int_81_174 bl_int_80_174 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c175
+ bl_int_81_175 bl_int_80_175 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c176
+ bl_int_81_176 bl_int_80_176 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c177
+ bl_int_81_177 bl_int_80_177 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c178
+ bl_int_81_178 bl_int_80_178 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c179
+ bl_int_81_179 bl_int_80_179 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c180
+ bl_int_81_180 bl_int_80_180 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c181
+ bl_int_81_181 bl_int_80_181 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c182
+ bl_int_81_182 bl_int_80_182 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r81_c183
+ bl_int_81_183 bl_int_80_183 wl_0_81 gnd
+ sram_rom_base_one_cell
Xbit_r82_c0
+ bl_int_82_0 bl_int_81_0 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c1
+ bl_int_82_1 bl_int_81_1 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c2
+ bl_int_82_2 bl_int_81_2 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c3
+ bl_int_82_3 bl_int_81_3 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c4
+ bl_int_82_4 bl_int_81_4 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c5
+ bl_int_82_5 bl_int_81_5 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c6
+ bl_int_82_6 bl_int_81_6 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c7
+ bl_int_82_7 bl_int_81_7 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c8
+ bl_int_82_8 bl_int_81_8 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c9
+ bl_int_82_9 bl_int_81_9 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c10
+ bl_int_82_10 bl_int_81_10 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c11
+ bl_int_82_11 bl_int_81_11 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c12
+ bl_int_82_12 bl_int_81_12 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c13
+ bl_int_82_13 bl_int_81_13 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c14
+ bl_int_82_14 bl_int_81_14 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c15
+ bl_int_82_15 bl_int_81_15 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c16
+ bl_int_82_16 bl_int_81_16 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c17
+ bl_int_82_17 bl_int_81_17 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c18
+ bl_int_82_18 bl_int_81_18 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c19
+ bl_int_82_19 bl_int_81_19 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c20
+ bl_int_82_20 bl_int_81_20 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c21
+ bl_int_82_21 bl_int_81_21 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c22
+ bl_int_82_22 bl_int_81_22 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c23
+ bl_int_82_23 bl_int_81_23 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c24
+ bl_int_82_24 bl_int_81_24 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c25
+ bl_int_82_25 bl_int_81_25 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c26
+ bl_int_82_26 bl_int_81_26 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c27
+ bl_int_82_27 bl_int_81_27 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c28
+ bl_int_82_28 bl_int_81_28 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c29
+ bl_int_82_29 bl_int_81_29 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c30
+ bl_int_82_30 bl_int_81_30 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c31
+ bl_int_82_31 bl_int_81_31 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c32
+ bl_int_82_32 bl_int_81_32 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c33
+ bl_int_82_33 bl_int_81_33 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c34
+ bl_int_82_34 bl_int_81_34 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c35
+ bl_int_82_35 bl_int_81_35 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c36
+ bl_int_82_36 bl_int_81_36 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c37
+ bl_int_82_37 bl_int_81_37 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c38
+ bl_int_82_38 bl_int_81_38 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c39
+ bl_int_82_39 bl_int_81_39 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c40
+ bl_int_82_40 bl_int_81_40 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c41
+ bl_int_82_41 bl_int_81_41 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c42
+ bl_int_82_42 bl_int_81_42 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c43
+ bl_int_82_43 bl_int_81_43 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c44
+ bl_int_82_44 bl_int_81_44 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c45
+ bl_int_82_45 bl_int_81_45 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c46
+ bl_int_82_46 bl_int_81_46 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c47
+ bl_int_82_47 bl_int_81_47 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c48
+ bl_int_82_48 bl_int_81_48 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c49
+ bl_int_82_49 bl_int_81_49 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c50
+ bl_int_82_50 bl_int_81_50 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c51
+ bl_int_82_51 bl_int_81_51 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c52
+ bl_int_82_52 bl_int_81_52 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c53
+ bl_int_82_53 bl_int_81_53 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c54
+ bl_int_82_54 bl_int_81_54 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c55
+ bl_int_82_55 bl_int_81_55 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c56
+ bl_int_82_56 bl_int_81_56 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c57
+ bl_int_82_57 bl_int_81_57 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c58
+ bl_int_82_58 bl_int_81_58 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c59
+ bl_int_82_59 bl_int_81_59 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c60
+ bl_int_82_60 bl_int_81_60 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c61
+ bl_int_82_61 bl_int_81_61 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c62
+ bl_int_82_62 bl_int_81_62 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c63
+ bl_int_82_63 bl_int_81_63 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c64
+ bl_int_82_64 bl_int_81_64 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c65
+ bl_int_82_65 bl_int_81_65 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c66
+ bl_int_82_66 bl_int_81_66 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c67
+ bl_int_82_67 bl_int_81_67 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c68
+ bl_int_82_68 bl_int_81_68 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c69
+ bl_int_82_69 bl_int_81_69 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c70
+ bl_int_82_70 bl_int_81_70 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c71
+ bl_int_82_71 bl_int_81_71 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c72
+ bl_int_82_72 bl_int_81_72 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c73
+ bl_int_82_73 bl_int_81_73 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c74
+ bl_int_82_74 bl_int_81_74 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c75
+ bl_int_82_75 bl_int_81_75 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c76
+ bl_int_82_76 bl_int_81_76 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c77
+ bl_int_82_77 bl_int_81_77 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c78
+ bl_int_82_78 bl_int_81_78 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c79
+ bl_int_82_79 bl_int_81_79 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c80
+ bl_int_82_80 bl_int_81_80 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c81
+ bl_int_82_81 bl_int_81_81 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c82
+ bl_int_82_82 bl_int_81_82 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c83
+ bl_int_82_83 bl_int_81_83 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c84
+ bl_int_82_84 bl_int_81_84 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c85
+ bl_int_82_85 bl_int_81_85 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c86
+ bl_int_82_86 bl_int_81_86 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c87
+ bl_int_82_87 bl_int_81_87 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c88
+ bl_int_82_88 bl_int_81_88 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c89
+ bl_int_82_89 bl_int_81_89 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c90
+ bl_int_82_90 bl_int_81_90 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c91
+ bl_int_82_91 bl_int_81_91 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c92
+ bl_int_82_92 bl_int_81_92 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c93
+ bl_int_82_93 bl_int_81_93 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c94
+ bl_int_82_94 bl_int_81_94 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c95
+ bl_int_82_95 bl_int_81_95 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c96
+ bl_int_82_96 bl_int_81_96 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c97
+ bl_int_82_97 bl_int_81_97 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c98
+ bl_int_82_98 bl_int_81_98 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c99
+ bl_int_82_99 bl_int_81_99 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c100
+ bl_int_82_100 bl_int_81_100 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c101
+ bl_int_82_101 bl_int_81_101 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c102
+ bl_int_82_102 bl_int_81_102 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c103
+ bl_int_82_103 bl_int_81_103 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c104
+ bl_int_82_104 bl_int_81_104 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c105
+ bl_int_82_105 bl_int_81_105 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c106
+ bl_int_82_106 bl_int_81_106 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c107
+ bl_int_82_107 bl_int_81_107 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c108
+ bl_int_82_108 bl_int_81_108 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c109
+ bl_int_82_109 bl_int_81_109 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c110
+ bl_int_82_110 bl_int_81_110 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c111
+ bl_int_82_111 bl_int_81_111 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c112
+ bl_int_82_112 bl_int_81_112 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c113
+ bl_int_82_113 bl_int_81_113 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c114
+ bl_int_82_114 bl_int_81_114 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c115
+ bl_int_82_115 bl_int_81_115 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c116
+ bl_int_82_116 bl_int_81_116 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c117
+ bl_int_82_117 bl_int_81_117 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c118
+ bl_int_82_118 bl_int_81_118 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c119
+ bl_int_82_119 bl_int_81_119 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c120
+ bl_int_82_120 bl_int_81_120 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c121
+ bl_int_82_121 bl_int_81_121 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c122
+ bl_int_82_122 bl_int_81_122 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c123
+ bl_int_82_123 bl_int_81_123 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c124
+ bl_int_82_124 bl_int_81_124 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c125
+ bl_int_82_125 bl_int_81_125 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c126
+ bl_int_82_126 bl_int_81_126 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c127
+ bl_int_82_127 bl_int_81_127 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c128
+ bl_int_82_128 bl_int_81_128 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c129
+ bl_int_82_129 bl_int_81_129 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c130
+ bl_int_82_130 bl_int_81_130 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c131
+ bl_int_82_131 bl_int_81_131 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c132
+ bl_int_82_132 bl_int_81_132 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c133
+ bl_int_82_133 bl_int_81_133 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c134
+ bl_int_82_134 bl_int_81_134 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c135
+ bl_int_82_135 bl_int_81_135 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c136
+ bl_int_82_136 bl_int_81_136 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c137
+ bl_int_82_137 bl_int_81_137 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c138
+ bl_int_82_138 bl_int_81_138 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c139
+ bl_int_82_139 bl_int_81_139 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c140
+ bl_int_82_140 bl_int_81_140 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c141
+ bl_int_82_141 bl_int_81_141 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c142
+ bl_int_82_142 bl_int_81_142 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c143
+ bl_int_82_143 bl_int_81_143 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c144
+ bl_int_82_144 bl_int_81_144 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c145
+ bl_int_82_145 bl_int_81_145 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c146
+ bl_int_82_146 bl_int_81_146 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c147
+ bl_int_82_147 bl_int_81_147 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c148
+ bl_int_82_148 bl_int_81_148 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c149
+ bl_int_82_149 bl_int_81_149 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c150
+ bl_int_82_150 bl_int_81_150 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c151
+ bl_int_82_151 bl_int_81_151 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c152
+ bl_int_82_152 bl_int_81_152 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c153
+ bl_int_82_153 bl_int_81_153 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c154
+ bl_int_82_154 bl_int_81_154 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c155
+ bl_int_82_155 bl_int_81_155 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c156
+ bl_int_82_156 bl_int_81_156 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c157
+ bl_int_82_157 bl_int_81_157 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c158
+ bl_int_82_158 bl_int_81_158 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c159
+ bl_int_82_159 bl_int_81_159 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c160
+ bl_int_82_160 bl_int_81_160 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c161
+ bl_int_82_161 bl_int_81_161 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c162
+ bl_int_82_162 bl_int_81_162 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c163
+ bl_int_82_163 bl_int_81_163 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c164
+ bl_int_82_164 bl_int_81_164 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c165
+ bl_int_82_165 bl_int_81_165 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c166
+ bl_int_82_166 bl_int_81_166 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c167
+ bl_int_82_167 bl_int_81_167 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c168
+ bl_int_82_168 bl_int_81_168 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c169
+ bl_int_82_169 bl_int_81_169 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c170
+ bl_int_82_170 bl_int_81_170 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c171
+ bl_int_82_171 bl_int_81_171 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c172
+ bl_int_82_172 bl_int_81_172 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c173
+ bl_int_82_173 bl_int_81_173 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c174
+ bl_int_82_174 bl_int_81_174 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c175
+ bl_int_82_175 bl_int_81_175 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c176
+ bl_int_82_176 bl_int_81_176 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c177
+ bl_int_82_177 bl_int_81_177 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c178
+ bl_int_82_178 bl_int_81_178 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c179
+ bl_int_82_179 bl_int_81_179 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c180
+ bl_int_82_180 bl_int_81_180 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c181
+ bl_int_82_181 bl_int_81_181 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c182
+ bl_int_82_182 bl_int_81_182 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r82_c183
+ bl_int_82_183 bl_int_81_183 wl_0_82 gnd
+ sram_rom_base_one_cell
Xbit_r83_c0
+ bl_int_83_0 bl_int_82_0 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c1
+ bl_int_83_1 bl_int_82_1 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c2
+ bl_int_83_2 bl_int_82_2 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c3
+ bl_int_83_3 bl_int_82_3 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c4
+ bl_int_83_4 bl_int_82_4 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c5
+ bl_int_83_5 bl_int_82_5 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c6
+ bl_int_83_6 bl_int_82_6 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c7
+ bl_int_83_7 bl_int_82_7 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c8
+ bl_int_83_8 bl_int_82_8 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c9
+ bl_int_83_9 bl_int_82_9 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c10
+ bl_int_83_10 bl_int_82_10 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c11
+ bl_int_83_11 bl_int_82_11 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c12
+ bl_int_83_12 bl_int_82_12 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c13
+ bl_int_83_13 bl_int_82_13 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c14
+ bl_int_83_14 bl_int_82_14 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c15
+ bl_int_83_15 bl_int_82_15 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c16
+ bl_int_83_16 bl_int_82_16 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c17
+ bl_int_83_17 bl_int_82_17 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c18
+ bl_int_83_18 bl_int_82_18 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c19
+ bl_int_83_19 bl_int_82_19 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c20
+ bl_int_83_20 bl_int_82_20 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c21
+ bl_int_83_21 bl_int_82_21 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c22
+ bl_int_83_22 bl_int_82_22 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c23
+ bl_int_83_23 bl_int_82_23 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c24
+ bl_int_83_24 bl_int_82_24 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c25
+ bl_int_83_25 bl_int_82_25 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c26
+ bl_int_83_26 bl_int_82_26 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c27
+ bl_int_83_27 bl_int_82_27 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c28
+ bl_int_83_28 bl_int_82_28 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c29
+ bl_int_83_29 bl_int_82_29 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c30
+ bl_int_83_30 bl_int_82_30 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c31
+ bl_int_83_31 bl_int_82_31 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c32
+ bl_int_83_32 bl_int_82_32 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c33
+ bl_int_83_33 bl_int_82_33 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c34
+ bl_int_83_34 bl_int_82_34 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c35
+ bl_int_83_35 bl_int_82_35 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c36
+ bl_int_83_36 bl_int_82_36 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c37
+ bl_int_83_37 bl_int_82_37 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c38
+ bl_int_83_38 bl_int_82_38 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c39
+ bl_int_83_39 bl_int_82_39 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c40
+ bl_int_83_40 bl_int_82_40 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c41
+ bl_int_83_41 bl_int_82_41 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c42
+ bl_int_83_42 bl_int_82_42 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c43
+ bl_int_83_43 bl_int_82_43 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c44
+ bl_int_83_44 bl_int_82_44 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c45
+ bl_int_83_45 bl_int_82_45 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c46
+ bl_int_83_46 bl_int_82_46 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c47
+ bl_int_83_47 bl_int_82_47 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c48
+ bl_int_83_48 bl_int_82_48 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c49
+ bl_int_83_49 bl_int_82_49 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c50
+ bl_int_83_50 bl_int_82_50 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c51
+ bl_int_83_51 bl_int_82_51 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c52
+ bl_int_83_52 bl_int_82_52 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c53
+ bl_int_83_53 bl_int_82_53 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c54
+ bl_int_83_54 bl_int_82_54 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c55
+ bl_int_83_55 bl_int_82_55 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c56
+ bl_int_83_56 bl_int_82_56 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c57
+ bl_int_83_57 bl_int_82_57 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c58
+ bl_int_83_58 bl_int_82_58 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c59
+ bl_int_83_59 bl_int_82_59 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c60
+ bl_int_83_60 bl_int_82_60 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c61
+ bl_int_83_61 bl_int_82_61 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c62
+ bl_int_83_62 bl_int_82_62 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c63
+ bl_int_83_63 bl_int_82_63 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c64
+ bl_int_83_64 bl_int_82_64 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c65
+ bl_int_83_65 bl_int_82_65 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c66
+ bl_int_83_66 bl_int_82_66 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c67
+ bl_int_83_67 bl_int_82_67 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c68
+ bl_int_83_68 bl_int_82_68 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c69
+ bl_int_83_69 bl_int_82_69 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c70
+ bl_int_83_70 bl_int_82_70 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c71
+ bl_int_83_71 bl_int_82_71 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c72
+ bl_int_83_72 bl_int_82_72 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c73
+ bl_int_83_73 bl_int_82_73 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c74
+ bl_int_83_74 bl_int_82_74 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c75
+ bl_int_83_75 bl_int_82_75 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c76
+ bl_int_83_76 bl_int_82_76 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c77
+ bl_int_83_77 bl_int_82_77 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c78
+ bl_int_83_78 bl_int_82_78 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c79
+ bl_int_83_79 bl_int_82_79 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c80
+ bl_int_83_80 bl_int_82_80 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c81
+ bl_int_83_81 bl_int_82_81 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c82
+ bl_int_83_82 bl_int_82_82 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c83
+ bl_int_83_83 bl_int_82_83 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c84
+ bl_int_83_84 bl_int_82_84 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c85
+ bl_int_83_85 bl_int_82_85 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c86
+ bl_int_83_86 bl_int_82_86 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c87
+ bl_int_83_87 bl_int_82_87 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c88
+ bl_int_83_88 bl_int_82_88 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c89
+ bl_int_83_89 bl_int_82_89 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c90
+ bl_int_83_90 bl_int_82_90 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c91
+ bl_int_83_91 bl_int_82_91 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c92
+ bl_int_83_92 bl_int_82_92 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c93
+ bl_int_83_93 bl_int_82_93 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c94
+ bl_int_83_94 bl_int_82_94 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c95
+ bl_int_83_95 bl_int_82_95 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c96
+ bl_int_83_96 bl_int_82_96 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c97
+ bl_int_83_97 bl_int_82_97 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c98
+ bl_int_83_98 bl_int_82_98 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c99
+ bl_int_83_99 bl_int_82_99 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c100
+ bl_int_83_100 bl_int_82_100 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c101
+ bl_int_83_101 bl_int_82_101 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c102
+ bl_int_83_102 bl_int_82_102 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c103
+ bl_int_83_103 bl_int_82_103 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c104
+ bl_int_83_104 bl_int_82_104 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c105
+ bl_int_83_105 bl_int_82_105 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c106
+ bl_int_83_106 bl_int_82_106 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c107
+ bl_int_83_107 bl_int_82_107 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c108
+ bl_int_83_108 bl_int_82_108 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c109
+ bl_int_83_109 bl_int_82_109 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c110
+ bl_int_83_110 bl_int_82_110 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c111
+ bl_int_83_111 bl_int_82_111 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c112
+ bl_int_83_112 bl_int_82_112 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c113
+ bl_int_83_113 bl_int_82_113 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c114
+ bl_int_83_114 bl_int_82_114 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c115
+ bl_int_83_115 bl_int_82_115 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c116
+ bl_int_83_116 bl_int_82_116 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c117
+ bl_int_83_117 bl_int_82_117 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c118
+ bl_int_83_118 bl_int_82_118 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c119
+ bl_int_83_119 bl_int_82_119 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c120
+ bl_int_83_120 bl_int_82_120 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c121
+ bl_int_83_121 bl_int_82_121 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c122
+ bl_int_83_122 bl_int_82_122 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c123
+ bl_int_83_123 bl_int_82_123 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c124
+ bl_int_83_124 bl_int_82_124 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c125
+ bl_int_83_125 bl_int_82_125 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c126
+ bl_int_83_126 bl_int_82_126 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c127
+ bl_int_83_127 bl_int_82_127 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c128
+ bl_int_83_128 bl_int_82_128 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c129
+ bl_int_83_129 bl_int_82_129 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c130
+ bl_int_83_130 bl_int_82_130 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c131
+ bl_int_83_131 bl_int_82_131 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c132
+ bl_int_83_132 bl_int_82_132 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c133
+ bl_int_83_133 bl_int_82_133 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c134
+ bl_int_83_134 bl_int_82_134 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c135
+ bl_int_83_135 bl_int_82_135 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c136
+ bl_int_83_136 bl_int_82_136 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c137
+ bl_int_83_137 bl_int_82_137 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c138
+ bl_int_83_138 bl_int_82_138 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c139
+ bl_int_83_139 bl_int_82_139 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c140
+ bl_int_83_140 bl_int_82_140 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c141
+ bl_int_83_141 bl_int_82_141 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c142
+ bl_int_83_142 bl_int_82_142 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c143
+ bl_int_83_143 bl_int_82_143 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c144
+ bl_int_83_144 bl_int_82_144 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c145
+ bl_int_83_145 bl_int_82_145 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c146
+ bl_int_83_146 bl_int_82_146 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c147
+ bl_int_83_147 bl_int_82_147 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c148
+ bl_int_83_148 bl_int_82_148 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c149
+ bl_int_83_149 bl_int_82_149 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c150
+ bl_int_83_150 bl_int_82_150 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c151
+ bl_int_83_151 bl_int_82_151 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c152
+ bl_int_83_152 bl_int_82_152 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c153
+ bl_int_83_153 bl_int_82_153 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c154
+ bl_int_83_154 bl_int_82_154 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c155
+ bl_int_83_155 bl_int_82_155 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c156
+ bl_int_83_156 bl_int_82_156 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c157
+ bl_int_83_157 bl_int_82_157 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c158
+ bl_int_83_158 bl_int_82_158 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c159
+ bl_int_83_159 bl_int_82_159 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c160
+ bl_int_83_160 bl_int_82_160 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c161
+ bl_int_83_161 bl_int_82_161 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c162
+ bl_int_83_162 bl_int_82_162 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c163
+ bl_int_83_163 bl_int_82_163 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c164
+ bl_int_83_164 bl_int_82_164 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c165
+ bl_int_83_165 bl_int_82_165 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c166
+ bl_int_83_166 bl_int_82_166 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c167
+ bl_int_83_167 bl_int_82_167 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c168
+ bl_int_83_168 bl_int_82_168 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c169
+ bl_int_83_169 bl_int_82_169 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c170
+ bl_int_83_170 bl_int_82_170 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c171
+ bl_int_83_171 bl_int_82_171 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c172
+ bl_int_83_172 bl_int_82_172 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c173
+ bl_int_83_173 bl_int_82_173 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c174
+ bl_int_83_174 bl_int_82_174 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c175
+ bl_int_83_175 bl_int_82_175 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c176
+ bl_int_83_176 bl_int_82_176 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c177
+ bl_int_83_177 bl_int_82_177 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c178
+ bl_int_83_178 bl_int_82_178 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c179
+ bl_int_83_179 bl_int_82_179 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c180
+ bl_int_83_180 bl_int_82_180 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c181
+ bl_int_83_181 bl_int_82_181 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c182
+ bl_int_83_182 bl_int_82_182 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r83_c183
+ bl_int_83_183 bl_int_82_183 wl_0_83 gnd
+ sram_rom_base_one_cell
Xbit_r84_c0
+ bl_int_84_0 bl_int_83_0 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c1
+ bl_int_84_1 bl_int_83_1 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c2
+ bl_int_84_2 bl_int_83_2 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c3
+ bl_int_84_3 bl_int_83_3 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c4
+ bl_int_84_4 bl_int_83_4 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c5
+ bl_int_84_5 bl_int_83_5 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c6
+ bl_int_84_6 bl_int_83_6 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c7
+ bl_int_84_7 bl_int_83_7 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c8
+ bl_int_84_8 bl_int_83_8 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c9
+ bl_int_84_9 bl_int_83_9 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c10
+ bl_int_84_10 bl_int_83_10 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c11
+ bl_int_84_11 bl_int_83_11 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c12
+ bl_int_84_12 bl_int_83_12 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c13
+ bl_int_84_13 bl_int_83_13 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c14
+ bl_int_84_14 bl_int_83_14 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c15
+ bl_int_84_15 bl_int_83_15 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c16
+ bl_int_84_16 bl_int_83_16 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c17
+ bl_int_84_17 bl_int_83_17 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c18
+ bl_int_84_18 bl_int_83_18 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c19
+ bl_int_84_19 bl_int_83_19 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c20
+ bl_int_84_20 bl_int_83_20 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c21
+ bl_int_84_21 bl_int_83_21 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c22
+ bl_int_84_22 bl_int_83_22 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c23
+ bl_int_84_23 bl_int_83_23 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c24
+ bl_int_84_24 bl_int_83_24 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c25
+ bl_int_84_25 bl_int_83_25 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c26
+ bl_int_84_26 bl_int_83_26 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c27
+ bl_int_84_27 bl_int_83_27 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c28
+ bl_int_84_28 bl_int_83_28 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c29
+ bl_int_84_29 bl_int_83_29 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c30
+ bl_int_84_30 bl_int_83_30 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c31
+ bl_int_84_31 bl_int_83_31 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c32
+ bl_int_84_32 bl_int_83_32 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c33
+ bl_int_84_33 bl_int_83_33 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c34
+ bl_int_84_34 bl_int_83_34 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c35
+ bl_int_84_35 bl_int_83_35 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c36
+ bl_int_84_36 bl_int_83_36 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c37
+ bl_int_84_37 bl_int_83_37 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c38
+ bl_int_84_38 bl_int_83_38 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c39
+ bl_int_84_39 bl_int_83_39 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c40
+ bl_int_84_40 bl_int_83_40 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c41
+ bl_int_84_41 bl_int_83_41 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c42
+ bl_int_84_42 bl_int_83_42 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c43
+ bl_int_84_43 bl_int_83_43 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c44
+ bl_int_84_44 bl_int_83_44 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c45
+ bl_int_84_45 bl_int_83_45 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c46
+ bl_int_84_46 bl_int_83_46 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c47
+ bl_int_84_47 bl_int_83_47 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c48
+ bl_int_84_48 bl_int_83_48 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c49
+ bl_int_84_49 bl_int_83_49 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c50
+ bl_int_84_50 bl_int_83_50 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c51
+ bl_int_84_51 bl_int_83_51 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c52
+ bl_int_84_52 bl_int_83_52 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c53
+ bl_int_84_53 bl_int_83_53 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c54
+ bl_int_84_54 bl_int_83_54 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c55
+ bl_int_84_55 bl_int_83_55 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c56
+ bl_int_84_56 bl_int_83_56 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c57
+ bl_int_84_57 bl_int_83_57 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c58
+ bl_int_84_58 bl_int_83_58 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c59
+ bl_int_84_59 bl_int_83_59 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c60
+ bl_int_84_60 bl_int_83_60 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c61
+ bl_int_84_61 bl_int_83_61 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c62
+ bl_int_84_62 bl_int_83_62 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c63
+ bl_int_84_63 bl_int_83_63 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c64
+ bl_int_84_64 bl_int_83_64 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c65
+ bl_int_84_65 bl_int_83_65 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c66
+ bl_int_84_66 bl_int_83_66 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c67
+ bl_int_84_67 bl_int_83_67 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c68
+ bl_int_84_68 bl_int_83_68 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c69
+ bl_int_84_69 bl_int_83_69 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c70
+ bl_int_84_70 bl_int_83_70 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c71
+ bl_int_84_71 bl_int_83_71 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c72
+ bl_int_84_72 bl_int_83_72 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c73
+ bl_int_84_73 bl_int_83_73 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c74
+ bl_int_84_74 bl_int_83_74 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c75
+ bl_int_84_75 bl_int_83_75 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c76
+ bl_int_84_76 bl_int_83_76 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c77
+ bl_int_84_77 bl_int_83_77 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c78
+ bl_int_84_78 bl_int_83_78 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c79
+ bl_int_84_79 bl_int_83_79 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c80
+ bl_int_84_80 bl_int_83_80 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c81
+ bl_int_84_81 bl_int_83_81 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c82
+ bl_int_84_82 bl_int_83_82 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c83
+ bl_int_84_83 bl_int_83_83 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c84
+ bl_int_84_84 bl_int_83_84 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c85
+ bl_int_84_85 bl_int_83_85 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c86
+ bl_int_84_86 bl_int_83_86 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c87
+ bl_int_84_87 bl_int_83_87 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c88
+ bl_int_84_88 bl_int_83_88 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c89
+ bl_int_84_89 bl_int_83_89 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c90
+ bl_int_84_90 bl_int_83_90 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c91
+ bl_int_84_91 bl_int_83_91 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c92
+ bl_int_84_92 bl_int_83_92 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c93
+ bl_int_84_93 bl_int_83_93 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c94
+ bl_int_84_94 bl_int_83_94 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c95
+ bl_int_84_95 bl_int_83_95 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c96
+ bl_int_84_96 bl_int_83_96 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c97
+ bl_int_84_97 bl_int_83_97 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c98
+ bl_int_84_98 bl_int_83_98 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c99
+ bl_int_84_99 bl_int_83_99 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c100
+ bl_int_84_100 bl_int_83_100 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c101
+ bl_int_84_101 bl_int_83_101 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c102
+ bl_int_84_102 bl_int_83_102 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c103
+ bl_int_84_103 bl_int_83_103 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c104
+ bl_int_84_104 bl_int_83_104 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c105
+ bl_int_84_105 bl_int_83_105 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c106
+ bl_int_84_106 bl_int_83_106 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c107
+ bl_int_84_107 bl_int_83_107 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c108
+ bl_int_84_108 bl_int_83_108 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c109
+ bl_int_84_109 bl_int_83_109 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c110
+ bl_int_84_110 bl_int_83_110 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c111
+ bl_int_84_111 bl_int_83_111 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c112
+ bl_int_84_112 bl_int_83_112 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c113
+ bl_int_84_113 bl_int_83_113 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c114
+ bl_int_84_114 bl_int_83_114 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c115
+ bl_int_84_115 bl_int_83_115 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c116
+ bl_int_84_116 bl_int_83_116 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c117
+ bl_int_84_117 bl_int_83_117 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c118
+ bl_int_84_118 bl_int_83_118 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c119
+ bl_int_84_119 bl_int_83_119 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c120
+ bl_int_84_120 bl_int_83_120 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c121
+ bl_int_84_121 bl_int_83_121 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c122
+ bl_int_84_122 bl_int_83_122 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c123
+ bl_int_84_123 bl_int_83_123 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c124
+ bl_int_84_124 bl_int_83_124 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c125
+ bl_int_84_125 bl_int_83_125 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c126
+ bl_int_84_126 bl_int_83_126 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c127
+ bl_int_84_127 bl_int_83_127 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c128
+ bl_int_84_128 bl_int_83_128 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c129
+ bl_int_84_129 bl_int_83_129 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c130
+ bl_int_84_130 bl_int_83_130 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c131
+ bl_int_84_131 bl_int_83_131 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c132
+ bl_int_84_132 bl_int_83_132 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c133
+ bl_int_84_133 bl_int_83_133 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c134
+ bl_int_84_134 bl_int_83_134 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c135
+ bl_int_84_135 bl_int_83_135 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c136
+ bl_int_84_136 bl_int_83_136 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c137
+ bl_int_84_137 bl_int_83_137 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c138
+ bl_int_84_138 bl_int_83_138 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c139
+ bl_int_84_139 bl_int_83_139 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c140
+ bl_int_84_140 bl_int_83_140 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c141
+ bl_int_84_141 bl_int_83_141 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c142
+ bl_int_84_142 bl_int_83_142 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c143
+ bl_int_84_143 bl_int_83_143 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c144
+ bl_int_84_144 bl_int_83_144 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c145
+ bl_int_84_145 bl_int_83_145 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c146
+ bl_int_84_146 bl_int_83_146 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c147
+ bl_int_84_147 bl_int_83_147 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c148
+ bl_int_84_148 bl_int_83_148 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c149
+ bl_int_84_149 bl_int_83_149 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c150
+ bl_int_84_150 bl_int_83_150 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c151
+ bl_int_84_151 bl_int_83_151 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c152
+ bl_int_84_152 bl_int_83_152 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c153
+ bl_int_84_153 bl_int_83_153 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c154
+ bl_int_84_154 bl_int_83_154 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c155
+ bl_int_84_155 bl_int_83_155 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c156
+ bl_int_84_156 bl_int_83_156 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c157
+ bl_int_84_157 bl_int_83_157 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c158
+ bl_int_84_158 bl_int_83_158 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c159
+ bl_int_84_159 bl_int_83_159 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c160
+ bl_int_84_160 bl_int_83_160 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c161
+ bl_int_84_161 bl_int_83_161 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c162
+ bl_int_84_162 bl_int_83_162 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c163
+ bl_int_84_163 bl_int_83_163 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c164
+ bl_int_84_164 bl_int_83_164 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c165
+ bl_int_84_165 bl_int_83_165 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c166
+ bl_int_84_166 bl_int_83_166 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c167
+ bl_int_84_167 bl_int_83_167 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c168
+ bl_int_84_168 bl_int_83_168 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c169
+ bl_int_84_169 bl_int_83_169 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c170
+ bl_int_84_170 bl_int_83_170 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c171
+ bl_int_84_171 bl_int_83_171 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c172
+ bl_int_84_172 bl_int_83_172 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c173
+ bl_int_84_173 bl_int_83_173 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c174
+ bl_int_84_174 bl_int_83_174 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c175
+ bl_int_84_175 bl_int_83_175 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c176
+ bl_int_84_176 bl_int_83_176 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c177
+ bl_int_84_177 bl_int_83_177 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c178
+ bl_int_84_178 bl_int_83_178 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c179
+ bl_int_84_179 bl_int_83_179 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c180
+ bl_int_84_180 bl_int_83_180 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c181
+ bl_int_84_181 bl_int_83_181 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c182
+ bl_int_84_182 bl_int_83_182 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r84_c183
+ bl_int_84_183 bl_int_83_183 wl_0_84 gnd
+ sram_rom_base_one_cell
Xbit_r85_c0
+ bl_int_85_0 bl_int_84_0 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c1
+ bl_int_85_1 bl_int_84_1 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c2
+ bl_int_85_2 bl_int_84_2 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c3
+ bl_int_85_3 bl_int_84_3 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c4
+ bl_int_85_4 bl_int_84_4 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c5
+ bl_int_85_5 bl_int_84_5 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c6
+ bl_int_85_6 bl_int_84_6 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c7
+ bl_int_85_7 bl_int_84_7 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c8
+ bl_int_85_8 bl_int_84_8 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c9
+ bl_int_85_9 bl_int_84_9 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c10
+ bl_int_85_10 bl_int_84_10 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c11
+ bl_int_85_11 bl_int_84_11 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c12
+ bl_int_85_12 bl_int_84_12 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c13
+ bl_int_85_13 bl_int_84_13 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c14
+ bl_int_85_14 bl_int_84_14 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c15
+ bl_int_85_15 bl_int_84_15 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c16
+ bl_int_85_16 bl_int_84_16 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c17
+ bl_int_85_17 bl_int_84_17 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c18
+ bl_int_85_18 bl_int_84_18 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c19
+ bl_int_85_19 bl_int_84_19 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c20
+ bl_int_85_20 bl_int_84_20 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c21
+ bl_int_85_21 bl_int_84_21 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c22
+ bl_int_85_22 bl_int_84_22 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c23
+ bl_int_85_23 bl_int_84_23 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c24
+ bl_int_85_24 bl_int_84_24 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c25
+ bl_int_85_25 bl_int_84_25 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c26
+ bl_int_85_26 bl_int_84_26 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c27
+ bl_int_85_27 bl_int_84_27 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c28
+ bl_int_85_28 bl_int_84_28 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c29
+ bl_int_85_29 bl_int_84_29 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c30
+ bl_int_85_30 bl_int_84_30 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c31
+ bl_int_85_31 bl_int_84_31 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c32
+ bl_int_85_32 bl_int_84_32 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c33
+ bl_int_85_33 bl_int_84_33 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c34
+ bl_int_85_34 bl_int_84_34 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c35
+ bl_int_85_35 bl_int_84_35 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c36
+ bl_int_85_36 bl_int_84_36 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c37
+ bl_int_85_37 bl_int_84_37 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c38
+ bl_int_85_38 bl_int_84_38 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c39
+ bl_int_85_39 bl_int_84_39 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c40
+ bl_int_85_40 bl_int_84_40 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c41
+ bl_int_85_41 bl_int_84_41 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c42
+ bl_int_85_42 bl_int_84_42 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c43
+ bl_int_85_43 bl_int_84_43 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c44
+ bl_int_85_44 bl_int_84_44 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c45
+ bl_int_85_45 bl_int_84_45 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c46
+ bl_int_85_46 bl_int_84_46 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c47
+ bl_int_85_47 bl_int_84_47 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c48
+ bl_int_85_48 bl_int_84_48 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c49
+ bl_int_85_49 bl_int_84_49 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c50
+ bl_int_85_50 bl_int_84_50 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c51
+ bl_int_85_51 bl_int_84_51 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c52
+ bl_int_85_52 bl_int_84_52 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c53
+ bl_int_85_53 bl_int_84_53 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c54
+ bl_int_85_54 bl_int_84_54 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c55
+ bl_int_85_55 bl_int_84_55 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c56
+ bl_int_85_56 bl_int_84_56 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c57
+ bl_int_85_57 bl_int_84_57 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c58
+ bl_int_85_58 bl_int_84_58 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c59
+ bl_int_85_59 bl_int_84_59 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c60
+ bl_int_85_60 bl_int_84_60 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c61
+ bl_int_85_61 bl_int_84_61 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c62
+ bl_int_85_62 bl_int_84_62 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c63
+ bl_int_85_63 bl_int_84_63 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c64
+ bl_int_85_64 bl_int_84_64 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c65
+ bl_int_85_65 bl_int_84_65 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c66
+ bl_int_85_66 bl_int_84_66 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c67
+ bl_int_85_67 bl_int_84_67 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c68
+ bl_int_85_68 bl_int_84_68 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c69
+ bl_int_85_69 bl_int_84_69 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c70
+ bl_int_85_70 bl_int_84_70 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c71
+ bl_int_85_71 bl_int_84_71 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c72
+ bl_int_85_72 bl_int_84_72 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c73
+ bl_int_85_73 bl_int_84_73 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c74
+ bl_int_85_74 bl_int_84_74 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c75
+ bl_int_85_75 bl_int_84_75 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c76
+ bl_int_85_76 bl_int_84_76 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c77
+ bl_int_85_77 bl_int_84_77 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c78
+ bl_int_85_78 bl_int_84_78 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c79
+ bl_int_85_79 bl_int_84_79 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c80
+ bl_int_85_80 bl_int_84_80 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c81
+ bl_int_85_81 bl_int_84_81 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c82
+ bl_int_85_82 bl_int_84_82 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c83
+ bl_int_85_83 bl_int_84_83 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c84
+ bl_int_85_84 bl_int_84_84 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c85
+ bl_int_85_85 bl_int_84_85 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c86
+ bl_int_85_86 bl_int_84_86 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c87
+ bl_int_85_87 bl_int_84_87 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c88
+ bl_int_85_88 bl_int_84_88 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c89
+ bl_int_85_89 bl_int_84_89 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c90
+ bl_int_85_90 bl_int_84_90 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c91
+ bl_int_85_91 bl_int_84_91 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c92
+ bl_int_85_92 bl_int_84_92 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c93
+ bl_int_85_93 bl_int_84_93 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c94
+ bl_int_85_94 bl_int_84_94 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c95
+ bl_int_85_95 bl_int_84_95 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c96
+ bl_int_85_96 bl_int_84_96 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c97
+ bl_int_85_97 bl_int_84_97 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c98
+ bl_int_85_98 bl_int_84_98 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c99
+ bl_int_85_99 bl_int_84_99 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c100
+ bl_int_85_100 bl_int_84_100 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c101
+ bl_int_85_101 bl_int_84_101 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c102
+ bl_int_85_102 bl_int_84_102 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c103
+ bl_int_85_103 bl_int_84_103 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c104
+ bl_int_85_104 bl_int_84_104 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c105
+ bl_int_85_105 bl_int_84_105 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c106
+ bl_int_85_106 bl_int_84_106 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c107
+ bl_int_85_107 bl_int_84_107 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c108
+ bl_int_85_108 bl_int_84_108 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c109
+ bl_int_85_109 bl_int_84_109 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c110
+ bl_int_85_110 bl_int_84_110 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c111
+ bl_int_85_111 bl_int_84_111 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c112
+ bl_int_85_112 bl_int_84_112 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c113
+ bl_int_85_113 bl_int_84_113 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c114
+ bl_int_85_114 bl_int_84_114 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c115
+ bl_int_85_115 bl_int_84_115 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c116
+ bl_int_85_116 bl_int_84_116 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c117
+ bl_int_85_117 bl_int_84_117 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c118
+ bl_int_85_118 bl_int_84_118 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c119
+ bl_int_85_119 bl_int_84_119 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c120
+ bl_int_85_120 bl_int_84_120 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c121
+ bl_int_85_121 bl_int_84_121 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c122
+ bl_int_85_122 bl_int_84_122 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c123
+ bl_int_85_123 bl_int_84_123 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c124
+ bl_int_85_124 bl_int_84_124 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c125
+ bl_int_85_125 bl_int_84_125 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c126
+ bl_int_85_126 bl_int_84_126 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c127
+ bl_int_85_127 bl_int_84_127 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c128
+ bl_int_85_128 bl_int_84_128 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c129
+ bl_int_85_129 bl_int_84_129 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c130
+ bl_int_85_130 bl_int_84_130 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c131
+ bl_int_85_131 bl_int_84_131 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c132
+ bl_int_85_132 bl_int_84_132 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c133
+ bl_int_85_133 bl_int_84_133 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c134
+ bl_int_85_134 bl_int_84_134 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c135
+ bl_int_85_135 bl_int_84_135 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c136
+ bl_int_85_136 bl_int_84_136 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c137
+ bl_int_85_137 bl_int_84_137 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c138
+ bl_int_85_138 bl_int_84_138 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c139
+ bl_int_85_139 bl_int_84_139 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c140
+ bl_int_85_140 bl_int_84_140 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c141
+ bl_int_85_141 bl_int_84_141 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c142
+ bl_int_85_142 bl_int_84_142 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c143
+ bl_int_85_143 bl_int_84_143 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c144
+ bl_int_85_144 bl_int_84_144 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c145
+ bl_int_85_145 bl_int_84_145 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c146
+ bl_int_85_146 bl_int_84_146 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c147
+ bl_int_85_147 bl_int_84_147 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c148
+ bl_int_85_148 bl_int_84_148 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c149
+ bl_int_85_149 bl_int_84_149 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c150
+ bl_int_85_150 bl_int_84_150 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c151
+ bl_int_85_151 bl_int_84_151 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c152
+ bl_int_85_152 bl_int_84_152 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c153
+ bl_int_85_153 bl_int_84_153 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c154
+ bl_int_85_154 bl_int_84_154 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c155
+ bl_int_85_155 bl_int_84_155 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c156
+ bl_int_85_156 bl_int_84_156 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c157
+ bl_int_85_157 bl_int_84_157 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c158
+ bl_int_85_158 bl_int_84_158 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c159
+ bl_int_85_159 bl_int_84_159 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c160
+ bl_int_85_160 bl_int_84_160 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c161
+ bl_int_85_161 bl_int_84_161 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c162
+ bl_int_85_162 bl_int_84_162 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c163
+ bl_int_85_163 bl_int_84_163 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c164
+ bl_int_85_164 bl_int_84_164 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c165
+ bl_int_85_165 bl_int_84_165 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c166
+ bl_int_85_166 bl_int_84_166 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c167
+ bl_int_85_167 bl_int_84_167 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c168
+ bl_int_85_168 bl_int_84_168 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c169
+ bl_int_85_169 bl_int_84_169 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c170
+ bl_int_85_170 bl_int_84_170 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c171
+ bl_int_85_171 bl_int_84_171 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c172
+ bl_int_85_172 bl_int_84_172 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c173
+ bl_int_85_173 bl_int_84_173 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c174
+ bl_int_85_174 bl_int_84_174 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c175
+ bl_int_85_175 bl_int_84_175 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c176
+ bl_int_85_176 bl_int_84_176 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c177
+ bl_int_85_177 bl_int_84_177 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c178
+ bl_int_85_178 bl_int_84_178 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c179
+ bl_int_85_179 bl_int_84_179 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c180
+ bl_int_85_180 bl_int_84_180 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c181
+ bl_int_85_181 bl_int_84_181 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c182
+ bl_int_85_182 bl_int_84_182 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r85_c183
+ bl_int_85_183 bl_int_84_183 wl_0_85 gnd
+ sram_rom_base_one_cell
Xbit_r86_c0
+ bl_int_86_0 bl_int_85_0 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c1
+ bl_int_86_1 bl_int_85_1 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c2
+ bl_int_86_2 bl_int_85_2 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c3
+ bl_int_86_3 bl_int_85_3 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c4
+ bl_int_86_4 bl_int_85_4 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c5
+ bl_int_86_5 bl_int_85_5 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c6
+ bl_int_86_6 bl_int_85_6 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c7
+ bl_int_86_7 bl_int_85_7 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c8
+ bl_int_86_8 bl_int_85_8 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c9
+ bl_int_86_9 bl_int_85_9 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c10
+ bl_int_86_10 bl_int_85_10 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c11
+ bl_int_86_11 bl_int_85_11 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c12
+ bl_int_86_12 bl_int_85_12 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c13
+ bl_int_86_13 bl_int_85_13 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c14
+ bl_int_86_14 bl_int_85_14 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c15
+ bl_int_86_15 bl_int_85_15 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c16
+ bl_int_86_16 bl_int_85_16 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c17
+ bl_int_86_17 bl_int_85_17 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c18
+ bl_int_86_18 bl_int_85_18 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c19
+ bl_int_86_19 bl_int_85_19 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c20
+ bl_int_86_20 bl_int_85_20 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c21
+ bl_int_86_21 bl_int_85_21 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c22
+ bl_int_86_22 bl_int_85_22 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c23
+ bl_int_86_23 bl_int_85_23 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c24
+ bl_int_86_24 bl_int_85_24 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c25
+ bl_int_86_25 bl_int_85_25 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c26
+ bl_int_86_26 bl_int_85_26 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c27
+ bl_int_86_27 bl_int_85_27 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c28
+ bl_int_86_28 bl_int_85_28 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c29
+ bl_int_86_29 bl_int_85_29 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c30
+ bl_int_86_30 bl_int_85_30 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c31
+ bl_int_86_31 bl_int_85_31 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c32
+ bl_int_86_32 bl_int_85_32 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c33
+ bl_int_86_33 bl_int_85_33 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c34
+ bl_int_86_34 bl_int_85_34 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c35
+ bl_int_86_35 bl_int_85_35 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c36
+ bl_int_86_36 bl_int_85_36 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c37
+ bl_int_86_37 bl_int_85_37 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c38
+ bl_int_86_38 bl_int_85_38 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c39
+ bl_int_86_39 bl_int_85_39 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c40
+ bl_int_86_40 bl_int_85_40 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c41
+ bl_int_86_41 bl_int_85_41 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c42
+ bl_int_86_42 bl_int_85_42 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c43
+ bl_int_86_43 bl_int_85_43 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c44
+ bl_int_86_44 bl_int_85_44 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c45
+ bl_int_86_45 bl_int_85_45 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c46
+ bl_int_86_46 bl_int_85_46 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c47
+ bl_int_86_47 bl_int_85_47 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c48
+ bl_int_86_48 bl_int_85_48 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c49
+ bl_int_86_49 bl_int_85_49 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c50
+ bl_int_86_50 bl_int_85_50 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c51
+ bl_int_86_51 bl_int_85_51 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c52
+ bl_int_86_52 bl_int_85_52 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c53
+ bl_int_86_53 bl_int_85_53 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c54
+ bl_int_86_54 bl_int_85_54 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c55
+ bl_int_86_55 bl_int_85_55 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c56
+ bl_int_86_56 bl_int_85_56 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c57
+ bl_int_86_57 bl_int_85_57 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c58
+ bl_int_86_58 bl_int_85_58 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c59
+ bl_int_86_59 bl_int_85_59 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c60
+ bl_int_86_60 bl_int_85_60 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c61
+ bl_int_86_61 bl_int_85_61 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c62
+ bl_int_86_62 bl_int_85_62 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c63
+ bl_int_86_63 bl_int_85_63 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c64
+ bl_int_86_64 bl_int_85_64 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c65
+ bl_int_86_65 bl_int_85_65 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c66
+ bl_int_86_66 bl_int_85_66 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c67
+ bl_int_86_67 bl_int_85_67 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c68
+ bl_int_86_68 bl_int_85_68 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c69
+ bl_int_86_69 bl_int_85_69 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c70
+ bl_int_86_70 bl_int_85_70 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c71
+ bl_int_86_71 bl_int_85_71 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c72
+ bl_int_86_72 bl_int_85_72 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c73
+ bl_int_86_73 bl_int_85_73 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c74
+ bl_int_86_74 bl_int_85_74 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c75
+ bl_int_86_75 bl_int_85_75 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c76
+ bl_int_86_76 bl_int_85_76 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c77
+ bl_int_86_77 bl_int_85_77 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c78
+ bl_int_86_78 bl_int_85_78 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c79
+ bl_int_86_79 bl_int_85_79 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c80
+ bl_int_86_80 bl_int_85_80 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c81
+ bl_int_86_81 bl_int_85_81 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c82
+ bl_int_86_82 bl_int_85_82 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c83
+ bl_int_86_83 bl_int_85_83 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c84
+ bl_int_86_84 bl_int_85_84 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c85
+ bl_int_86_85 bl_int_85_85 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c86
+ bl_int_86_86 bl_int_85_86 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c87
+ bl_int_86_87 bl_int_85_87 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c88
+ bl_int_86_88 bl_int_85_88 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c89
+ bl_int_86_89 bl_int_85_89 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c90
+ bl_int_86_90 bl_int_85_90 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c91
+ bl_int_86_91 bl_int_85_91 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c92
+ bl_int_86_92 bl_int_85_92 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c93
+ bl_int_86_93 bl_int_85_93 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c94
+ bl_int_86_94 bl_int_85_94 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c95
+ bl_int_86_95 bl_int_85_95 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c96
+ bl_int_86_96 bl_int_85_96 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c97
+ bl_int_86_97 bl_int_85_97 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c98
+ bl_int_86_98 bl_int_85_98 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c99
+ bl_int_86_99 bl_int_85_99 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c100
+ bl_int_86_100 bl_int_85_100 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c101
+ bl_int_86_101 bl_int_85_101 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c102
+ bl_int_86_102 bl_int_85_102 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c103
+ bl_int_86_103 bl_int_85_103 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c104
+ bl_int_86_104 bl_int_85_104 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c105
+ bl_int_86_105 bl_int_85_105 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c106
+ bl_int_86_106 bl_int_85_106 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c107
+ bl_int_86_107 bl_int_85_107 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c108
+ bl_int_86_108 bl_int_85_108 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c109
+ bl_int_86_109 bl_int_85_109 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c110
+ bl_int_86_110 bl_int_85_110 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c111
+ bl_int_86_111 bl_int_85_111 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c112
+ bl_int_86_112 bl_int_85_112 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c113
+ bl_int_86_113 bl_int_85_113 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c114
+ bl_int_86_114 bl_int_85_114 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c115
+ bl_int_86_115 bl_int_85_115 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c116
+ bl_int_86_116 bl_int_85_116 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c117
+ bl_int_86_117 bl_int_85_117 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c118
+ bl_int_86_118 bl_int_85_118 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c119
+ bl_int_86_119 bl_int_85_119 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c120
+ bl_int_86_120 bl_int_85_120 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c121
+ bl_int_86_121 bl_int_85_121 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c122
+ bl_int_86_122 bl_int_85_122 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c123
+ bl_int_86_123 bl_int_85_123 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c124
+ bl_int_86_124 bl_int_85_124 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c125
+ bl_int_86_125 bl_int_85_125 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c126
+ bl_int_86_126 bl_int_85_126 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c127
+ bl_int_86_127 bl_int_85_127 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c128
+ bl_int_86_128 bl_int_85_128 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c129
+ bl_int_86_129 bl_int_85_129 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c130
+ bl_int_86_130 bl_int_85_130 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c131
+ bl_int_86_131 bl_int_85_131 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c132
+ bl_int_86_132 bl_int_85_132 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c133
+ bl_int_86_133 bl_int_85_133 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c134
+ bl_int_86_134 bl_int_85_134 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c135
+ bl_int_86_135 bl_int_85_135 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c136
+ bl_int_86_136 bl_int_85_136 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c137
+ bl_int_86_137 bl_int_85_137 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c138
+ bl_int_86_138 bl_int_85_138 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c139
+ bl_int_86_139 bl_int_85_139 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c140
+ bl_int_86_140 bl_int_85_140 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c141
+ bl_int_86_141 bl_int_85_141 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c142
+ bl_int_86_142 bl_int_85_142 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c143
+ bl_int_86_143 bl_int_85_143 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c144
+ bl_int_86_144 bl_int_85_144 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c145
+ bl_int_86_145 bl_int_85_145 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c146
+ bl_int_86_146 bl_int_85_146 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c147
+ bl_int_86_147 bl_int_85_147 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c148
+ bl_int_86_148 bl_int_85_148 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c149
+ bl_int_86_149 bl_int_85_149 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c150
+ bl_int_86_150 bl_int_85_150 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c151
+ bl_int_86_151 bl_int_85_151 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c152
+ bl_int_86_152 bl_int_85_152 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c153
+ bl_int_86_153 bl_int_85_153 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c154
+ bl_int_86_154 bl_int_85_154 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c155
+ bl_int_86_155 bl_int_85_155 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c156
+ bl_int_86_156 bl_int_85_156 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c157
+ bl_int_86_157 bl_int_85_157 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c158
+ bl_int_86_158 bl_int_85_158 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c159
+ bl_int_86_159 bl_int_85_159 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c160
+ bl_int_86_160 bl_int_85_160 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c161
+ bl_int_86_161 bl_int_85_161 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c162
+ bl_int_86_162 bl_int_85_162 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c163
+ bl_int_86_163 bl_int_85_163 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c164
+ bl_int_86_164 bl_int_85_164 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c165
+ bl_int_86_165 bl_int_85_165 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c166
+ bl_int_86_166 bl_int_85_166 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c167
+ bl_int_86_167 bl_int_85_167 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c168
+ bl_int_86_168 bl_int_85_168 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c169
+ bl_int_86_169 bl_int_85_169 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c170
+ bl_int_86_170 bl_int_85_170 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c171
+ bl_int_86_171 bl_int_85_171 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c172
+ bl_int_86_172 bl_int_85_172 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c173
+ bl_int_86_173 bl_int_85_173 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c174
+ bl_int_86_174 bl_int_85_174 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c175
+ bl_int_86_175 bl_int_85_175 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c176
+ bl_int_86_176 bl_int_85_176 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c177
+ bl_int_86_177 bl_int_85_177 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c178
+ bl_int_86_178 bl_int_85_178 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c179
+ bl_int_86_179 bl_int_85_179 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c180
+ bl_int_86_180 bl_int_85_180 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c181
+ bl_int_86_181 bl_int_85_181 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c182
+ bl_int_86_182 bl_int_85_182 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r86_c183
+ bl_int_86_183 bl_int_85_183 wl_0_86 gnd
+ sram_rom_base_one_cell
Xbit_r87_c0
+ bl_int_87_0 bl_int_86_0 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c1
+ bl_int_87_1 bl_int_86_1 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c2
+ bl_int_87_2 bl_int_86_2 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c3
+ bl_int_87_3 bl_int_86_3 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c4
+ bl_int_87_4 bl_int_86_4 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c5
+ bl_int_87_5 bl_int_86_5 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c6
+ bl_int_87_6 bl_int_86_6 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c7
+ bl_int_87_7 bl_int_86_7 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c8
+ bl_int_87_8 bl_int_86_8 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c9
+ bl_int_87_9 bl_int_86_9 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c10
+ bl_int_87_10 bl_int_86_10 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c11
+ bl_int_87_11 bl_int_86_11 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c12
+ bl_int_87_12 bl_int_86_12 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c13
+ bl_int_87_13 bl_int_86_13 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c14
+ bl_int_87_14 bl_int_86_14 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c15
+ bl_int_86_15 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c16
+ bl_int_86_16 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c17
+ bl_int_86_17 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c18
+ bl_int_86_18 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c19
+ bl_int_86_19 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c20
+ bl_int_86_20 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c21
+ bl_int_86_21 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c22
+ bl_int_86_22 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c23
+ bl_int_87_23 bl_int_86_23 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c24
+ bl_int_87_24 bl_int_86_24 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c25
+ bl_int_87_25 bl_int_86_25 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c26
+ bl_int_87_26 bl_int_86_26 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c27
+ bl_int_87_27 bl_int_86_27 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c28
+ bl_int_87_28 bl_int_86_28 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c29
+ bl_int_87_29 bl_int_86_29 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c30
+ bl_int_87_30 bl_int_86_30 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c31
+ bl_int_87_31 bl_int_86_31 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c32
+ bl_int_87_32 bl_int_86_32 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c33
+ bl_int_87_33 bl_int_86_33 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c34
+ bl_int_87_34 bl_int_86_34 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c35
+ bl_int_87_35 bl_int_86_35 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c36
+ bl_int_87_36 bl_int_86_36 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c37
+ bl_int_87_37 bl_int_86_37 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c38
+ bl_int_86_38 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c39
+ bl_int_86_39 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c40
+ bl_int_86_40 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c41
+ bl_int_86_41 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c42
+ bl_int_86_42 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c43
+ bl_int_86_43 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c44
+ bl_int_86_44 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c45
+ bl_int_86_45 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c46
+ bl_int_87_46 bl_int_86_46 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c47
+ bl_int_87_47 bl_int_86_47 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c48
+ bl_int_87_48 bl_int_86_48 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c49
+ bl_int_87_49 bl_int_86_49 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c50
+ bl_int_87_50 bl_int_86_50 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c51
+ bl_int_87_51 bl_int_86_51 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c52
+ bl_int_87_52 bl_int_86_52 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c53
+ bl_int_87_53 bl_int_86_53 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c54
+ bl_int_87_54 bl_int_86_54 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c55
+ bl_int_87_55 bl_int_86_55 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c56
+ bl_int_87_56 bl_int_86_56 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c57
+ bl_int_87_57 bl_int_86_57 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c58
+ bl_int_87_58 bl_int_86_58 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c59
+ bl_int_87_59 bl_int_86_59 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c60
+ bl_int_87_60 bl_int_86_60 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c61
+ bl_int_86_61 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c62
+ bl_int_86_62 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c63
+ bl_int_86_63 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c64
+ bl_int_86_64 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c65
+ bl_int_86_65 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c66
+ bl_int_86_66 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c67
+ bl_int_86_67 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c68
+ bl_int_86_68 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c69
+ bl_int_87_69 bl_int_86_69 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c70
+ bl_int_87_70 bl_int_86_70 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c71
+ bl_int_87_71 bl_int_86_71 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c72
+ bl_int_87_72 bl_int_86_72 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c73
+ bl_int_87_73 bl_int_86_73 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c74
+ bl_int_87_74 bl_int_86_74 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c75
+ bl_int_87_75 bl_int_86_75 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c76
+ bl_int_87_76 bl_int_86_76 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c77
+ bl_int_87_77 bl_int_86_77 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c78
+ bl_int_87_78 bl_int_86_78 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c79
+ bl_int_87_79 bl_int_86_79 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c80
+ bl_int_87_80 bl_int_86_80 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c81
+ bl_int_87_81 bl_int_86_81 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c82
+ bl_int_87_82 bl_int_86_82 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c83
+ bl_int_87_83 bl_int_86_83 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c84
+ bl_int_86_84 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c85
+ bl_int_86_85 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c86
+ bl_int_86_86 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c87
+ bl_int_86_87 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c88
+ bl_int_86_88 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c89
+ bl_int_86_89 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c90
+ bl_int_86_90 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c91
+ bl_int_86_91 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c92
+ bl_int_87_92 bl_int_86_92 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c93
+ bl_int_87_93 bl_int_86_93 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c94
+ bl_int_87_94 bl_int_86_94 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c95
+ bl_int_87_95 bl_int_86_95 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c96
+ bl_int_87_96 bl_int_86_96 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c97
+ bl_int_87_97 bl_int_86_97 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c98
+ bl_int_87_98 bl_int_86_98 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c99
+ bl_int_87_99 bl_int_86_99 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c100
+ bl_int_87_100 bl_int_86_100 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c101
+ bl_int_87_101 bl_int_86_101 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c102
+ bl_int_87_102 bl_int_86_102 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c103
+ bl_int_87_103 bl_int_86_103 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c104
+ bl_int_87_104 bl_int_86_104 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c105
+ bl_int_87_105 bl_int_86_105 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c106
+ bl_int_87_106 bl_int_86_106 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c107
+ bl_int_86_107 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c108
+ bl_int_86_108 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c109
+ bl_int_86_109 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c110
+ bl_int_86_110 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c111
+ bl_int_86_111 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c112
+ bl_int_86_112 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c113
+ bl_int_86_113 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c114
+ bl_int_86_114 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c115
+ bl_int_87_115 bl_int_86_115 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c116
+ bl_int_87_116 bl_int_86_116 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c117
+ bl_int_87_117 bl_int_86_117 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c118
+ bl_int_87_118 bl_int_86_118 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c119
+ bl_int_87_119 bl_int_86_119 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c120
+ bl_int_87_120 bl_int_86_120 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c121
+ bl_int_87_121 bl_int_86_121 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c122
+ bl_int_87_122 bl_int_86_122 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c123
+ bl_int_87_123 bl_int_86_123 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c124
+ bl_int_87_124 bl_int_86_124 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c125
+ bl_int_87_125 bl_int_86_125 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c126
+ bl_int_87_126 bl_int_86_126 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c127
+ bl_int_87_127 bl_int_86_127 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c128
+ bl_int_87_128 bl_int_86_128 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c129
+ bl_int_87_129 bl_int_86_129 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c130
+ bl_int_86_130 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c131
+ bl_int_86_131 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c132
+ bl_int_86_132 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c133
+ bl_int_86_133 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c134
+ bl_int_86_134 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c135
+ bl_int_86_135 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c136
+ bl_int_86_136 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c137
+ bl_int_86_137 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c138
+ bl_int_87_138 bl_int_86_138 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c139
+ bl_int_87_139 bl_int_86_139 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c140
+ bl_int_87_140 bl_int_86_140 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c141
+ bl_int_87_141 bl_int_86_141 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c142
+ bl_int_87_142 bl_int_86_142 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c143
+ bl_int_87_143 bl_int_86_143 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c144
+ bl_int_87_144 bl_int_86_144 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c145
+ bl_int_87_145 bl_int_86_145 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c146
+ bl_int_87_146 bl_int_86_146 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c147
+ bl_int_87_147 bl_int_86_147 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c148
+ bl_int_87_148 bl_int_86_148 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c149
+ bl_int_87_149 bl_int_86_149 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c150
+ bl_int_87_150 bl_int_86_150 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c151
+ bl_int_87_151 bl_int_86_151 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c152
+ bl_int_87_152 bl_int_86_152 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c153
+ bl_int_86_153 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c154
+ bl_int_86_154 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c155
+ bl_int_86_155 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c156
+ bl_int_86_156 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c157
+ bl_int_86_157 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c158
+ bl_int_86_158 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c159
+ bl_int_86_159 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c160
+ bl_int_86_160 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c161
+ bl_int_87_161 bl_int_86_161 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c162
+ bl_int_87_162 bl_int_86_162 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c163
+ bl_int_87_163 bl_int_86_163 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c164
+ bl_int_87_164 bl_int_86_164 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c165
+ bl_int_87_165 bl_int_86_165 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c166
+ bl_int_87_166 bl_int_86_166 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c167
+ bl_int_87_167 bl_int_86_167 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c168
+ bl_int_87_168 bl_int_86_168 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c169
+ bl_int_87_169 bl_int_86_169 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c170
+ bl_int_87_170 bl_int_86_170 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c171
+ bl_int_87_171 bl_int_86_171 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c172
+ bl_int_87_172 bl_int_86_172 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c173
+ bl_int_87_173 bl_int_86_173 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c174
+ bl_int_87_174 bl_int_86_174 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c175
+ bl_int_87_175 bl_int_86_175 wl_0_87 gnd
+ sram_rom_base_one_cell
Xbit_r87_c176
+ bl_int_86_176 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c177
+ bl_int_86_177 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c178
+ bl_int_86_178 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c179
+ bl_int_86_179 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c180
+ bl_int_86_180 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c181
+ bl_int_86_181 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c182
+ bl_int_86_182 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r87_c183
+ bl_int_86_183 wl_0_87 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c0
+ bl_int_87_0 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c1
+ bl_int_87_1 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c2
+ bl_int_87_2 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c3
+ bl_int_87_3 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c4
+ bl_int_87_4 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c5
+ bl_int_87_5 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c6
+ bl_int_87_6 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c7
+ bl_int_87_7 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c8
+ bl_int_88_8 bl_int_87_8 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c9
+ bl_int_88_9 bl_int_87_9 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c10
+ bl_int_88_10 bl_int_87_10 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c11
+ bl_int_88_11 bl_int_87_11 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c12
+ bl_int_88_12 bl_int_87_12 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c13
+ bl_int_88_13 bl_int_87_13 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c14
+ bl_int_88_14 bl_int_87_14 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c15
+ bl_int_88_15 bl_int_86_15 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c16
+ bl_int_88_16 bl_int_86_16 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c17
+ bl_int_88_17 bl_int_86_17 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c18
+ bl_int_88_18 bl_int_86_18 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c19
+ bl_int_88_19 bl_int_86_19 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c20
+ bl_int_88_20 bl_int_86_20 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c21
+ bl_int_88_21 bl_int_86_21 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c22
+ bl_int_88_22 bl_int_86_22 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c23
+ bl_int_87_23 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c24
+ bl_int_87_24 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c25
+ bl_int_87_25 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c26
+ bl_int_87_26 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c27
+ bl_int_87_27 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c28
+ bl_int_87_28 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c29
+ bl_int_87_29 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c30
+ bl_int_87_30 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c31
+ bl_int_88_31 bl_int_87_31 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c32
+ bl_int_88_32 bl_int_87_32 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c33
+ bl_int_88_33 bl_int_87_33 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c34
+ bl_int_88_34 bl_int_87_34 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c35
+ bl_int_88_35 bl_int_87_35 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c36
+ bl_int_88_36 bl_int_87_36 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c37
+ bl_int_88_37 bl_int_87_37 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c38
+ bl_int_88_38 bl_int_86_38 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c39
+ bl_int_88_39 bl_int_86_39 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c40
+ bl_int_88_40 bl_int_86_40 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c41
+ bl_int_88_41 bl_int_86_41 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c42
+ bl_int_88_42 bl_int_86_42 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c43
+ bl_int_88_43 bl_int_86_43 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c44
+ bl_int_88_44 bl_int_86_44 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c45
+ bl_int_88_45 bl_int_86_45 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c46
+ bl_int_87_46 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c47
+ bl_int_87_47 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c48
+ bl_int_87_48 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c49
+ bl_int_87_49 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c50
+ bl_int_87_50 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c51
+ bl_int_87_51 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c52
+ bl_int_87_52 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c53
+ bl_int_87_53 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c54
+ bl_int_88_54 bl_int_87_54 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c55
+ bl_int_88_55 bl_int_87_55 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c56
+ bl_int_88_56 bl_int_87_56 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c57
+ bl_int_88_57 bl_int_87_57 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c58
+ bl_int_88_58 bl_int_87_58 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c59
+ bl_int_88_59 bl_int_87_59 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c60
+ bl_int_88_60 bl_int_87_60 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c61
+ bl_int_88_61 bl_int_86_61 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c62
+ bl_int_88_62 bl_int_86_62 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c63
+ bl_int_88_63 bl_int_86_63 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c64
+ bl_int_88_64 bl_int_86_64 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c65
+ bl_int_88_65 bl_int_86_65 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c66
+ bl_int_88_66 bl_int_86_66 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c67
+ bl_int_88_67 bl_int_86_67 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c68
+ bl_int_88_68 bl_int_86_68 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c69
+ bl_int_87_69 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c70
+ bl_int_87_70 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c71
+ bl_int_87_71 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c72
+ bl_int_87_72 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c73
+ bl_int_87_73 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c74
+ bl_int_87_74 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c75
+ bl_int_87_75 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c76
+ bl_int_87_76 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c77
+ bl_int_88_77 bl_int_87_77 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c78
+ bl_int_88_78 bl_int_87_78 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c79
+ bl_int_88_79 bl_int_87_79 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c80
+ bl_int_88_80 bl_int_87_80 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c81
+ bl_int_88_81 bl_int_87_81 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c82
+ bl_int_88_82 bl_int_87_82 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c83
+ bl_int_88_83 bl_int_87_83 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c84
+ bl_int_88_84 bl_int_86_84 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c85
+ bl_int_88_85 bl_int_86_85 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c86
+ bl_int_88_86 bl_int_86_86 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c87
+ bl_int_88_87 bl_int_86_87 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c88
+ bl_int_88_88 bl_int_86_88 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c89
+ bl_int_88_89 bl_int_86_89 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c90
+ bl_int_88_90 bl_int_86_90 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c91
+ bl_int_88_91 bl_int_86_91 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c92
+ bl_int_87_92 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c93
+ bl_int_87_93 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c94
+ bl_int_87_94 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c95
+ bl_int_87_95 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c96
+ bl_int_87_96 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c97
+ bl_int_87_97 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c98
+ bl_int_87_98 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c99
+ bl_int_87_99 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c100
+ bl_int_88_100 bl_int_87_100 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c101
+ bl_int_88_101 bl_int_87_101 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c102
+ bl_int_88_102 bl_int_87_102 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c103
+ bl_int_88_103 bl_int_87_103 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c104
+ bl_int_88_104 bl_int_87_104 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c105
+ bl_int_88_105 bl_int_87_105 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c106
+ bl_int_88_106 bl_int_87_106 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c107
+ bl_int_88_107 bl_int_86_107 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c108
+ bl_int_88_108 bl_int_86_108 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c109
+ bl_int_88_109 bl_int_86_109 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c110
+ bl_int_88_110 bl_int_86_110 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c111
+ bl_int_88_111 bl_int_86_111 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c112
+ bl_int_88_112 bl_int_86_112 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c113
+ bl_int_88_113 bl_int_86_113 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c114
+ bl_int_88_114 bl_int_86_114 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c115
+ bl_int_87_115 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c116
+ bl_int_87_116 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c117
+ bl_int_87_117 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c118
+ bl_int_87_118 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c119
+ bl_int_87_119 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c120
+ bl_int_87_120 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c121
+ bl_int_87_121 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c122
+ bl_int_87_122 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c123
+ bl_int_88_123 bl_int_87_123 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c124
+ bl_int_88_124 bl_int_87_124 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c125
+ bl_int_88_125 bl_int_87_125 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c126
+ bl_int_88_126 bl_int_87_126 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c127
+ bl_int_88_127 bl_int_87_127 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c128
+ bl_int_88_128 bl_int_87_128 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c129
+ bl_int_88_129 bl_int_87_129 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c130
+ bl_int_88_130 bl_int_86_130 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c131
+ bl_int_88_131 bl_int_86_131 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c132
+ bl_int_88_132 bl_int_86_132 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c133
+ bl_int_88_133 bl_int_86_133 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c134
+ bl_int_88_134 bl_int_86_134 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c135
+ bl_int_88_135 bl_int_86_135 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c136
+ bl_int_88_136 bl_int_86_136 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c137
+ bl_int_88_137 bl_int_86_137 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c138
+ bl_int_87_138 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c139
+ bl_int_87_139 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c140
+ bl_int_87_140 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c141
+ bl_int_87_141 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c142
+ bl_int_87_142 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c143
+ bl_int_87_143 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c144
+ bl_int_87_144 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c145
+ bl_int_87_145 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c146
+ bl_int_88_146 bl_int_87_146 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c147
+ bl_int_88_147 bl_int_87_147 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c148
+ bl_int_88_148 bl_int_87_148 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c149
+ bl_int_88_149 bl_int_87_149 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c150
+ bl_int_88_150 bl_int_87_150 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c151
+ bl_int_88_151 bl_int_87_151 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c152
+ bl_int_88_152 bl_int_87_152 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c153
+ bl_int_88_153 bl_int_86_153 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c154
+ bl_int_88_154 bl_int_86_154 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c155
+ bl_int_88_155 bl_int_86_155 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c156
+ bl_int_88_156 bl_int_86_156 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c157
+ bl_int_88_157 bl_int_86_157 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c158
+ bl_int_88_158 bl_int_86_158 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c159
+ bl_int_88_159 bl_int_86_159 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c160
+ bl_int_88_160 bl_int_86_160 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c161
+ bl_int_87_161 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c162
+ bl_int_87_162 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c163
+ bl_int_87_163 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c164
+ bl_int_87_164 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c165
+ bl_int_87_165 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c166
+ bl_int_87_166 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c167
+ bl_int_87_167 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c168
+ bl_int_87_168 wl_0_88 gnd
+ sram_rom_base_zero_cell
Xbit_r88_c169
+ bl_int_88_169 bl_int_87_169 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c170
+ bl_int_88_170 bl_int_87_170 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c171
+ bl_int_88_171 bl_int_87_171 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c172
+ bl_int_88_172 bl_int_87_172 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c173
+ bl_int_88_173 bl_int_87_173 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c174
+ bl_int_88_174 bl_int_87_174 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c175
+ bl_int_88_175 bl_int_87_175 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c176
+ bl_int_88_176 bl_int_86_176 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c177
+ bl_int_88_177 bl_int_86_177 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c178
+ bl_int_88_178 bl_int_86_178 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c179
+ bl_int_88_179 bl_int_86_179 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c180
+ bl_int_88_180 bl_int_86_180 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c181
+ bl_int_88_181 bl_int_86_181 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c182
+ bl_int_88_182 bl_int_86_182 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r88_c183
+ bl_int_88_183 bl_int_86_183 wl_0_88 gnd
+ sram_rom_base_one_cell
Xbit_r89_c0
+ gnd bl_int_87_0 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c1
+ gnd bl_int_87_1 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c2
+ gnd bl_int_87_2 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c3
+ gnd bl_int_87_3 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c4
+ gnd bl_int_87_4 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c5
+ gnd bl_int_87_5 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c6
+ gnd bl_int_87_6 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c7
+ gnd bl_int_87_7 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c8
+ gnd bl_int_88_8 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c9
+ gnd bl_int_88_9 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c10
+ gnd bl_int_88_10 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c11
+ gnd bl_int_88_11 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c12
+ gnd bl_int_88_12 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c13
+ gnd bl_int_88_13 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c14
+ gnd bl_int_88_14 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c15
+ gnd bl_int_88_15 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c16
+ gnd bl_int_88_16 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c17
+ gnd bl_int_88_17 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c18
+ gnd bl_int_88_18 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c19
+ gnd bl_int_88_19 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c20
+ gnd bl_int_88_20 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c21
+ gnd bl_int_88_21 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c22
+ gnd bl_int_88_22 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c23
+ gnd bl_int_87_23 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c24
+ gnd bl_int_87_24 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c25
+ gnd bl_int_87_25 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c26
+ gnd bl_int_87_26 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c27
+ gnd bl_int_87_27 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c28
+ gnd bl_int_87_28 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c29
+ gnd bl_int_87_29 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c30
+ gnd bl_int_87_30 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c31
+ gnd bl_int_88_31 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c32
+ gnd bl_int_88_32 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c33
+ gnd bl_int_88_33 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c34
+ gnd bl_int_88_34 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c35
+ gnd bl_int_88_35 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c36
+ gnd bl_int_88_36 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c37
+ gnd bl_int_88_37 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c38
+ gnd bl_int_88_38 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c39
+ gnd bl_int_88_39 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c40
+ gnd bl_int_88_40 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c41
+ gnd bl_int_88_41 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c42
+ gnd bl_int_88_42 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c43
+ gnd bl_int_88_43 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c44
+ gnd bl_int_88_44 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c45
+ gnd bl_int_88_45 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c46
+ gnd bl_int_87_46 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c47
+ gnd bl_int_87_47 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c48
+ gnd bl_int_87_48 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c49
+ gnd bl_int_87_49 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c50
+ gnd bl_int_87_50 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c51
+ gnd bl_int_87_51 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c52
+ gnd bl_int_87_52 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c53
+ gnd bl_int_87_53 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c54
+ gnd bl_int_88_54 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c55
+ gnd bl_int_88_55 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c56
+ gnd bl_int_88_56 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c57
+ gnd bl_int_88_57 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c58
+ gnd bl_int_88_58 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c59
+ gnd bl_int_88_59 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c60
+ gnd bl_int_88_60 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c61
+ gnd bl_int_88_61 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c62
+ gnd bl_int_88_62 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c63
+ gnd bl_int_88_63 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c64
+ gnd bl_int_88_64 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c65
+ gnd bl_int_88_65 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c66
+ gnd bl_int_88_66 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c67
+ gnd bl_int_88_67 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c68
+ gnd bl_int_88_68 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c69
+ gnd bl_int_87_69 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c70
+ gnd bl_int_87_70 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c71
+ gnd bl_int_87_71 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c72
+ gnd bl_int_87_72 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c73
+ gnd bl_int_87_73 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c74
+ gnd bl_int_87_74 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c75
+ gnd bl_int_87_75 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c76
+ gnd bl_int_87_76 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c77
+ gnd bl_int_88_77 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c78
+ gnd bl_int_88_78 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c79
+ gnd bl_int_88_79 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c80
+ gnd bl_int_88_80 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c81
+ gnd bl_int_88_81 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c82
+ gnd bl_int_88_82 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c83
+ gnd bl_int_88_83 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c84
+ gnd bl_int_88_84 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c85
+ gnd bl_int_88_85 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c86
+ gnd bl_int_88_86 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c87
+ gnd bl_int_88_87 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c88
+ gnd bl_int_88_88 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c89
+ gnd bl_int_88_89 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c90
+ gnd bl_int_88_90 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c91
+ gnd bl_int_88_91 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c92
+ gnd bl_int_87_92 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c93
+ gnd bl_int_87_93 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c94
+ gnd bl_int_87_94 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c95
+ gnd bl_int_87_95 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c96
+ gnd bl_int_87_96 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c97
+ gnd bl_int_87_97 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c98
+ gnd bl_int_87_98 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c99
+ gnd bl_int_87_99 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c100
+ gnd bl_int_88_100 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c101
+ gnd bl_int_88_101 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c102
+ gnd bl_int_88_102 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c103
+ gnd bl_int_88_103 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c104
+ gnd bl_int_88_104 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c105
+ gnd bl_int_88_105 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c106
+ gnd bl_int_88_106 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c107
+ gnd bl_int_88_107 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c108
+ gnd bl_int_88_108 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c109
+ gnd bl_int_88_109 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c110
+ gnd bl_int_88_110 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c111
+ gnd bl_int_88_111 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c112
+ gnd bl_int_88_112 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c113
+ gnd bl_int_88_113 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c114
+ gnd bl_int_88_114 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c115
+ gnd bl_int_87_115 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c116
+ gnd bl_int_87_116 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c117
+ gnd bl_int_87_117 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c118
+ gnd bl_int_87_118 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c119
+ gnd bl_int_87_119 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c120
+ gnd bl_int_87_120 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c121
+ gnd bl_int_87_121 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c122
+ gnd bl_int_87_122 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c123
+ gnd bl_int_88_123 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c124
+ gnd bl_int_88_124 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c125
+ gnd bl_int_88_125 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c126
+ gnd bl_int_88_126 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c127
+ gnd bl_int_88_127 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c128
+ gnd bl_int_88_128 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c129
+ gnd bl_int_88_129 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c130
+ gnd bl_int_88_130 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c131
+ gnd bl_int_88_131 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c132
+ gnd bl_int_88_132 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c133
+ gnd bl_int_88_133 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c134
+ gnd bl_int_88_134 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c135
+ gnd bl_int_88_135 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c136
+ gnd bl_int_88_136 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c137
+ gnd bl_int_88_137 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c138
+ gnd bl_int_87_138 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c139
+ gnd bl_int_87_139 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c140
+ gnd bl_int_87_140 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c141
+ gnd bl_int_87_141 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c142
+ gnd bl_int_87_142 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c143
+ gnd bl_int_87_143 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c144
+ gnd bl_int_87_144 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c145
+ gnd bl_int_87_145 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c146
+ gnd bl_int_88_146 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c147
+ gnd bl_int_88_147 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c148
+ gnd bl_int_88_148 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c149
+ gnd bl_int_88_149 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c150
+ gnd bl_int_88_150 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c151
+ gnd bl_int_88_151 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c152
+ gnd bl_int_88_152 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c153
+ gnd bl_int_88_153 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c154
+ gnd bl_int_88_154 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c155
+ gnd bl_int_88_155 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c156
+ gnd bl_int_88_156 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c157
+ gnd bl_int_88_157 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c158
+ gnd bl_int_88_158 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c159
+ gnd bl_int_88_159 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c160
+ gnd bl_int_88_160 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c161
+ gnd bl_int_87_161 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c162
+ gnd bl_int_87_162 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c163
+ gnd bl_int_87_163 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c164
+ gnd bl_int_87_164 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c165
+ gnd bl_int_87_165 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c166
+ gnd bl_int_87_166 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c167
+ gnd bl_int_87_167 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c168
+ gnd bl_int_87_168 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c169
+ gnd bl_int_88_169 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c170
+ gnd bl_int_88_170 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c171
+ gnd bl_int_88_171 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c172
+ gnd bl_int_88_172 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c173
+ gnd bl_int_88_173 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c174
+ gnd bl_int_88_174 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c175
+ gnd bl_int_88_175 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c176
+ gnd bl_int_88_176 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c177
+ gnd bl_int_88_177 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c178
+ gnd bl_int_88_178 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c179
+ gnd bl_int_88_179 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c180
+ gnd bl_int_88_180 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c181
+ gnd bl_int_88_181 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c182
+ gnd bl_int_88_182 precharge gnd
+ sram_rom_base_one_cell
Xbit_r89_c183
+ gnd bl_int_88_183 precharge gnd
+ sram_rom_base_one_cell
Xbitcell_array_precharge
+ bl_0_0 bl_0_1 bl_0_2 bl_0_3 bl_0_4 bl_0_5 bl_0_6 bl_0_7 bl_0_8 bl_0_9
+ bl_0_10 bl_0_11 bl_0_12 bl_0_13 bl_0_14 bl_0_15 bl_0_16 bl_0_17
+ bl_0_18 bl_0_19 bl_0_20 bl_0_21 bl_0_22 bl_0_23 bl_0_24 bl_0_25
+ bl_0_26 bl_0_27 bl_0_28 bl_0_29 bl_0_30 bl_0_31 bl_0_32 bl_0_33
+ bl_0_34 bl_0_35 bl_0_36 bl_0_37 bl_0_38 bl_0_39 bl_0_40 bl_0_41
+ bl_0_42 bl_0_43 bl_0_44 bl_0_45 bl_0_46 bl_0_47 bl_0_48 bl_0_49
+ bl_0_50 bl_0_51 bl_0_52 bl_0_53 bl_0_54 bl_0_55 bl_0_56 bl_0_57
+ bl_0_58 bl_0_59 bl_0_60 bl_0_61 bl_0_62 bl_0_63 bl_0_64 bl_0_65
+ bl_0_66 bl_0_67 bl_0_68 bl_0_69 bl_0_70 bl_0_71 bl_0_72 bl_0_73
+ bl_0_74 bl_0_75 bl_0_76 bl_0_77 bl_0_78 bl_0_79 bl_0_80 bl_0_81
+ bl_0_82 bl_0_83 bl_0_84 bl_0_85 bl_0_86 bl_0_87 bl_0_88 bl_0_89
+ bl_0_90 bl_0_91 bl_0_92 bl_0_93 bl_0_94 bl_0_95 bl_0_96 bl_0_97
+ bl_0_98 bl_0_99 bl_0_100 bl_0_101 bl_0_102 bl_0_103 bl_0_104 bl_0_105
+ bl_0_106 bl_0_107 bl_0_108 bl_0_109 bl_0_110 bl_0_111 bl_0_112
+ bl_0_113 bl_0_114 bl_0_115 bl_0_116 bl_0_117 bl_0_118 bl_0_119
+ bl_0_120 bl_0_121 bl_0_122 bl_0_123 bl_0_124 bl_0_125 bl_0_126
+ bl_0_127 bl_0_128 bl_0_129 bl_0_130 bl_0_131 bl_0_132 bl_0_133
+ bl_0_134 bl_0_135 bl_0_136 bl_0_137 bl_0_138 bl_0_139 bl_0_140
+ bl_0_141 bl_0_142 bl_0_143 bl_0_144 bl_0_145 bl_0_146 bl_0_147
+ bl_0_148 bl_0_149 bl_0_150 bl_0_151 bl_0_152 bl_0_153 bl_0_154
+ bl_0_155 bl_0_156 bl_0_157 bl_0_158 bl_0_159 bl_0_160 bl_0_161
+ bl_0_162 bl_0_163 bl_0_164 bl_0_165 bl_0_166 bl_0_167 bl_0_168
+ bl_0_169 bl_0_170 bl_0_171 bl_0_172 bl_0_173 bl_0_174 bl_0_175
+ bl_0_176 bl_0_177 bl_0_178 bl_0_179 bl_0_180 bl_0_181 bl_0_182
+ bl_0_183 precharge vdd
+ sram_rom_precharge_array
.ENDS sram_rom_base_array

.SUBCKT sram_rom_base_bank
+ clk CS addr_0 addr_1 addr_2 addr_3 addr_4 addr_5 addr_6 addr_7 addr_8
+ addr_9 addr_10 addr_11 rom_out_0 rom_out_1 rom_out_2 rom_out_3
+ rom_out_4 rom_out_5 rom_out_6 rom_out_7 vdd gnd
* INPUT : clk 
* INPUT : CS 
* INPUT : addr_0 
* INPUT : addr_1 
* INPUT : addr_2 
* INPUT : addr_3 
* INPUT : addr_4 
* INPUT : addr_5 
* INPUT : addr_6 
* INPUT : addr_7 
* INPUT : addr_8 
* INPUT : addr_9 
* INPUT : addr_10 
* INPUT : addr_11 
* OUTPUT: rom_out_0 
* OUTPUT: rom_out_1 
* OUTPUT: rom_out_2 
* OUTPUT: rom_out_3 
* OUTPUT: rom_out_4 
* OUTPUT: rom_out_5 
* OUTPUT: rom_out_6 
* OUTPUT: rom_out_7 
* POWER : vdd 
* GROUND: gnd 
Xrom_bit_array
+ bl_0 bl_1 bl_2 bl_3 bl_4 bl_5 bl_6 bl_7 bl_8 bl_9 bl_10 bl_11 bl_12
+ bl_13 bl_14 bl_15 bl_16 bl_17 bl_18 bl_19 bl_20 bl_21 bl_22 bl_23
+ bl_24 bl_25 bl_26 bl_27 bl_28 bl_29 bl_30 bl_31 bl_32 bl_33 bl_34
+ bl_35 bl_36 bl_37 bl_38 bl_39 bl_40 bl_41 bl_42 bl_43 bl_44 bl_45
+ bl_46 bl_47 bl_48 bl_49 bl_50 bl_51 bl_52 bl_53 bl_54 bl_55 bl_56
+ bl_57 bl_58 bl_59 bl_60 bl_61 bl_62 bl_63 bl_64 bl_65 bl_66 bl_67
+ bl_68 bl_69 bl_70 bl_71 bl_72 bl_73 bl_74 bl_75 bl_76 bl_77 bl_78
+ bl_79 bl_80 bl_81 bl_82 bl_83 bl_84 bl_85 bl_86 bl_87 bl_88 bl_89
+ bl_90 bl_91 bl_92 bl_93 bl_94 bl_95 bl_96 bl_97 bl_98 bl_99 bl_100
+ bl_101 bl_102 bl_103 bl_104 bl_105 bl_106 bl_107 bl_108 bl_109 bl_110
+ bl_111 bl_112 bl_113 bl_114 bl_115 bl_116 bl_117 bl_118 bl_119 bl_120
+ bl_121 bl_122 bl_123 bl_124 bl_125 bl_126 bl_127 bl_128 bl_129 bl_130
+ bl_131 bl_132 bl_133 bl_134 bl_135 bl_136 bl_137 bl_138 bl_139 bl_140
+ bl_141 bl_142 bl_143 bl_144 bl_145 bl_146 bl_147 bl_148 bl_149 bl_150
+ bl_151 bl_152 bl_153 bl_154 bl_155 bl_156 bl_157 bl_158 bl_159 bl_160
+ bl_161 bl_162 bl_163 bl_164 bl_165 bl_166 bl_167 bl_168 bl_169 bl_170
+ bl_171 bl_172 bl_173 bl_174 bl_175 bl_176 bl_177 bl_178 bl_179 bl_180
+ bl_181 bl_182 bl_183 wl_0 wl_1 wl_2 wl_3 wl_4 wl_5 wl_6 wl_7 wl_8 wl_9
+ wl_10 wl_11 wl_12 wl_13 wl_14 wl_15 wl_16 wl_17 wl_18 wl_19 wl_20
+ wl_21 wl_22 wl_23 wl_24 wl_25 wl_26 wl_27 wl_28 wl_29 wl_30 wl_31
+ wl_32 wl_33 wl_34 wl_35 wl_36 wl_37 wl_38 wl_39 wl_40 wl_41 wl_42
+ wl_43 wl_44 wl_45 wl_46 wl_47 wl_48 wl_49 wl_50 wl_51 wl_52 wl_53
+ wl_54 wl_55 wl_56 wl_57 wl_58 wl_59 wl_60 wl_61 wl_62 wl_63 wl_64
+ wl_65 wl_66 wl_67 wl_68 wl_69 wl_70 wl_71 wl_72 wl_73 wl_74 wl_75
+ wl_76 wl_77 wl_78 wl_79 wl_80 wl_81 wl_82 wl_83 wl_84 wl_85 wl_86
+ wl_87 wl_88 precharge vdd gnd
+ sram_rom_base_array
Xrom_row_decoder
+ addr_5 addr_6 addr_7 addr_8 addr_9 addr_10 addr_11 wl_0 wl_1 wl_2 wl_3
+ wl_4 wl_5 wl_6 wl_7 wl_8 wl_9 wl_10 wl_11 wl_12 wl_13 wl_14 wl_15
+ wl_16 wl_17 wl_18 wl_19 wl_20 wl_21 wl_22 wl_23 wl_24 wl_25 wl_26
+ wl_27 wl_28 wl_29 wl_30 wl_31 wl_32 wl_33 wl_34 wl_35 wl_36 wl_37
+ wl_38 wl_39 wl_40 wl_41 wl_42 wl_43 wl_44 wl_45 wl_46 wl_47 wl_48
+ wl_49 wl_50 wl_51 wl_52 wl_53 wl_54 wl_55 wl_56 wl_57 wl_58 wl_59
+ wl_60 wl_61 wl_62 wl_63 wl_64 wl_65 wl_66 wl_67 wl_68 wl_69 wl_70
+ wl_71 wl_72 wl_73 wl_74 wl_75 wl_76 wl_77 wl_78 wl_79 wl_80 wl_81
+ wl_82 wl_83 wl_84 wl_85 wl_86 wl_87 wl_88 clk_int clk_int vdd gnd
+ sram_rom_row_decode
Xrom_control
+ clk CS precharge clk_int vdd gnd
+ sram_rom_control_logic
Xrom_column_mux
+ bl_b_0 bl_b_1 bl_b_2 bl_b_3 bl_b_4 bl_b_5 bl_b_6 bl_b_7 bl_b_8 bl_b_9
+ bl_b_10 bl_b_11 bl_b_12 bl_b_13 bl_b_14 bl_b_15 bl_b_16 bl_b_17
+ bl_b_18 bl_b_19 bl_b_20 bl_b_21 bl_b_22 bl_b_23 bl_b_24 bl_b_25
+ bl_b_26 bl_b_27 bl_b_28 bl_b_29 bl_b_30 bl_b_31 bl_b_32 bl_b_33
+ bl_b_34 bl_b_35 bl_b_36 bl_b_37 bl_b_38 bl_b_39 bl_b_40 bl_b_41
+ bl_b_42 bl_b_43 bl_b_44 bl_b_45 bl_b_46 bl_b_47 bl_b_48 bl_b_49
+ bl_b_50 bl_b_51 bl_b_52 bl_b_53 bl_b_54 bl_b_55 bl_b_56 bl_b_57
+ bl_b_58 bl_b_59 bl_b_60 bl_b_61 bl_b_62 bl_b_63 bl_b_64 bl_b_65
+ bl_b_66 bl_b_67 bl_b_68 bl_b_69 bl_b_70 bl_b_71 bl_b_72 bl_b_73
+ bl_b_74 bl_b_75 bl_b_76 bl_b_77 bl_b_78 bl_b_79 bl_b_80 bl_b_81
+ bl_b_82 bl_b_83 bl_b_84 bl_b_85 bl_b_86 bl_b_87 bl_b_88 bl_b_89
+ bl_b_90 bl_b_91 bl_b_92 bl_b_93 bl_b_94 bl_b_95 bl_b_96 bl_b_97
+ bl_b_98 bl_b_99 bl_b_100 bl_b_101 bl_b_102 bl_b_103 bl_b_104 bl_b_105
+ bl_b_106 bl_b_107 bl_b_108 bl_b_109 bl_b_110 bl_b_111 bl_b_112
+ bl_b_113 bl_b_114 bl_b_115 bl_b_116 bl_b_117 bl_b_118 bl_b_119
+ bl_b_120 bl_b_121 bl_b_122 bl_b_123 bl_b_124 bl_b_125 bl_b_126
+ bl_b_127 bl_b_128 bl_b_129 bl_b_130 bl_b_131 bl_b_132 bl_b_133
+ bl_b_134 bl_b_135 bl_b_136 bl_b_137 bl_b_138 bl_b_139 bl_b_140
+ bl_b_141 bl_b_142 bl_b_143 bl_b_144 bl_b_145 bl_b_146 bl_b_147
+ bl_b_148 bl_b_149 bl_b_150 bl_b_151 bl_b_152 bl_b_153 bl_b_154
+ bl_b_155 bl_b_156 bl_b_157 bl_b_158 bl_b_159 bl_b_160 bl_b_161
+ bl_b_162 bl_b_163 bl_b_164 bl_b_165 bl_b_166 bl_b_167 bl_b_168
+ bl_b_169 bl_b_170 bl_b_171 bl_b_172 bl_b_173 bl_b_174 bl_b_175
+ bl_b_176 bl_b_177 bl_b_178 bl_b_179 bl_b_180 bl_b_181 bl_b_182
+ bl_b_183 word_sel_0 word_sel_1 word_sel_2 word_sel_3 word_sel_4
+ word_sel_5 word_sel_6 word_sel_7 word_sel_8 word_sel_9 word_sel_10
+ word_sel_11 word_sel_12 word_sel_13 word_sel_14 word_sel_15
+ word_sel_16 word_sel_17 word_sel_18 word_sel_19 word_sel_20
+ word_sel_21 word_sel_22 rom_out_prebuf_0 rom_out_prebuf_1
+ rom_out_prebuf_2 rom_out_prebuf_3 rom_out_prebuf_4 rom_out_prebuf_5
+ rom_out_prebuf_6 rom_out_prebuf_7 gnd
+ sram_rom_column_mux_array
Xrom_column_decoder
+ addr_0 addr_1 addr_2 addr_3 addr_4 word_sel_0 word_sel_1 word_sel_2
+ word_sel_3 word_sel_4 word_sel_5 word_sel_6 word_sel_7 word_sel_8
+ word_sel_9 word_sel_10 word_sel_11 word_sel_12 word_sel_13 word_sel_14
+ word_sel_15 word_sel_16 word_sel_17 word_sel_18 word_sel_19
+ word_sel_20 word_sel_21 word_sel_22 precharge precharge vdd gnd
+ sram_rom_column_decode
Xrom_bitline_inverter
+ bl_0 bl_1 bl_2 bl_3 bl_4 bl_5 bl_6 bl_7 bl_8 bl_9 bl_10 bl_11 bl_12
+ bl_13 bl_14 bl_15 bl_16 bl_17 bl_18 bl_19 bl_20 bl_21 bl_22 bl_23
+ bl_24 bl_25 bl_26 bl_27 bl_28 bl_29 bl_30 bl_31 bl_32 bl_33 bl_34
+ bl_35 bl_36 bl_37 bl_38 bl_39 bl_40 bl_41 bl_42 bl_43 bl_44 bl_45
+ bl_46 bl_47 bl_48 bl_49 bl_50 bl_51 bl_52 bl_53 bl_54 bl_55 bl_56
+ bl_57 bl_58 bl_59 bl_60 bl_61 bl_62 bl_63 bl_64 bl_65 bl_66 bl_67
+ bl_68 bl_69 bl_70 bl_71 bl_72 bl_73 bl_74 bl_75 bl_76 bl_77 bl_78
+ bl_79 bl_80 bl_81 bl_82 bl_83 bl_84 bl_85 bl_86 bl_87 bl_88 bl_89
+ bl_90 bl_91 bl_92 bl_93 bl_94 bl_95 bl_96 bl_97 bl_98 bl_99 bl_100
+ bl_101 bl_102 bl_103 bl_104 bl_105 bl_106 bl_107 bl_108 bl_109 bl_110
+ bl_111 bl_112 bl_113 bl_114 bl_115 bl_116 bl_117 bl_118 bl_119 bl_120
+ bl_121 bl_122 bl_123 bl_124 bl_125 bl_126 bl_127 bl_128 bl_129 bl_130
+ bl_131 bl_132 bl_133 bl_134 bl_135 bl_136 bl_137 bl_138 bl_139 bl_140
+ bl_141 bl_142 bl_143 bl_144 bl_145 bl_146 bl_147 bl_148 bl_149 bl_150
+ bl_151 bl_152 bl_153 bl_154 bl_155 bl_156 bl_157 bl_158 bl_159 bl_160
+ bl_161 bl_162 bl_163 bl_164 bl_165 bl_166 bl_167 bl_168 bl_169 bl_170
+ bl_171 bl_172 bl_173 bl_174 bl_175 bl_176 bl_177 bl_178 bl_179 bl_180
+ bl_181 bl_182 bl_183 bl_b_0 bl_b_1 bl_b_2 bl_b_3 bl_b_4 bl_b_5 bl_b_6
+ bl_b_7 bl_b_8 bl_b_9 bl_b_10 bl_b_11 bl_b_12 bl_b_13 bl_b_14 bl_b_15
+ bl_b_16 bl_b_17 bl_b_18 bl_b_19 bl_b_20 bl_b_21 bl_b_22 bl_b_23
+ bl_b_24 bl_b_25 bl_b_26 bl_b_27 bl_b_28 bl_b_29 bl_b_30 bl_b_31
+ bl_b_32 bl_b_33 bl_b_34 bl_b_35 bl_b_36 bl_b_37 bl_b_38 bl_b_39
+ bl_b_40 bl_b_41 bl_b_42 bl_b_43 bl_b_44 bl_b_45 bl_b_46 bl_b_47
+ bl_b_48 bl_b_49 bl_b_50 bl_b_51 bl_b_52 bl_b_53 bl_b_54 bl_b_55
+ bl_b_56 bl_b_57 bl_b_58 bl_b_59 bl_b_60 bl_b_61 bl_b_62 bl_b_63
+ bl_b_64 bl_b_65 bl_b_66 bl_b_67 bl_b_68 bl_b_69 bl_b_70 bl_b_71
+ bl_b_72 bl_b_73 bl_b_74 bl_b_75 bl_b_76 bl_b_77 bl_b_78 bl_b_79
+ bl_b_80 bl_b_81 bl_b_82 bl_b_83 bl_b_84 bl_b_85 bl_b_86 bl_b_87
+ bl_b_88 bl_b_89 bl_b_90 bl_b_91 bl_b_92 bl_b_93 bl_b_94 bl_b_95
+ bl_b_96 bl_b_97 bl_b_98 bl_b_99 bl_b_100 bl_b_101 bl_b_102 bl_b_103
+ bl_b_104 bl_b_105 bl_b_106 bl_b_107 bl_b_108 bl_b_109 bl_b_110
+ bl_b_111 bl_b_112 bl_b_113 bl_b_114 bl_b_115 bl_b_116 bl_b_117
+ bl_b_118 bl_b_119 bl_b_120 bl_b_121 bl_b_122 bl_b_123 bl_b_124
+ bl_b_125 bl_b_126 bl_b_127 bl_b_128 bl_b_129 bl_b_130 bl_b_131
+ bl_b_132 bl_b_133 bl_b_134 bl_b_135 bl_b_136 bl_b_137 bl_b_138
+ bl_b_139 bl_b_140 bl_b_141 bl_b_142 bl_b_143 bl_b_144 bl_b_145
+ bl_b_146 bl_b_147 bl_b_148 bl_b_149 bl_b_150 bl_b_151 bl_b_152
+ bl_b_153 bl_b_154 bl_b_155 bl_b_156 bl_b_157 bl_b_158 bl_b_159
+ bl_b_160 bl_b_161 bl_b_162 bl_b_163 bl_b_164 bl_b_165 bl_b_166
+ bl_b_167 bl_b_168 bl_b_169 bl_b_170 bl_b_171 bl_b_172 bl_b_173
+ bl_b_174 bl_b_175 bl_b_176 bl_b_177 bl_b_178 bl_b_179 bl_b_180
+ bl_b_181 bl_b_182 bl_b_183 vdd gnd
+ sram_rom_bitline_inverter
Xrom_output_inverter
+ rom_out_prebuf_0 rom_out_prebuf_1 rom_out_prebuf_2 rom_out_prebuf_3
+ rom_out_prebuf_4 rom_out_prebuf_5 rom_out_prebuf_6 rom_out_prebuf_7
+ rom_out_0 rom_out_1 rom_out_2 rom_out_3 rom_out_4 rom_out_5 rom_out_6
+ rom_out_7 vdd gnd
+ sram_rom_output_buffer
.ENDS sram_rom_base_bank
